
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;
USE std.env.finish;

ENTITY random_tb IS
END random_tb;

ARCHITECTURE randomtb OF random_tb IS
	CONSTANT CLOCK_PERIOD : TIME := 100 ns;
	SIGNAL tb_done : STD_LOGIC;
	SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
	SIGNAL tb_rst : STD_LOGIC := '0';
	SIGNAL tb_start : STD_LOGIC := '0';
	SIGNAL tb_clk : STD_LOGIC := '0';
	SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL enable_wire : STD_LOGIC;
	SIGNAL mem_we : STD_LOGIC;
	SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL tb_w : STD_LOGIC;

	CONSTANT SCENARIOLENGTH : INTEGER := 405951;
	CONSTANT N_EVENTS : INTEGER := 10000;
	SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)		:= "010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)	:= "010011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000001111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000001111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000011111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000101111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000011111111111111111000000000000000000000001111111111100000000000000000000000111111111111111000000000000000000000001111111111111111100000000000000000000100000111111111111111111000000000000000000000000111111111111111110000000000000000000010011111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000010000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000001000011111111111111111100000000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000010111111111111111110000000000000000000010001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111000000000000000000001000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111110000000000000000000000000111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100001111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000010001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111100000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000010000011111111111111111000000000000000000000111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111100000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000001001111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000010111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000011111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000100111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000010000111111111111111110000000000000000000010111111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000100001111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000000111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000101111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111110000000000000000000001111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111000000000000000000001000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000010001111111111111111110000000000000000000010000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000001011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010001111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000010001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010000011111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000011111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111110000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001001111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000010011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111000000000000000000000011111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111110000000000000000000000111111111111111111000000000000000000000001111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000100001111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001000111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010000011111111111111110000000000000000000010000011111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000100001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000010000011111111111111111100000000000000000000101111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000001000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001000011111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000010000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010001111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000100000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000001001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000010111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000010001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000111111111111111100000000000000000000000000111111111111111110000000000000000000010111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001011111111111111110000000000000000000010011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000010011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000001011111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000010111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000001011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000001111111111111111100000000000000000000100000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000001000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000010000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000010000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000100001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000001111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000010011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111110000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111100000000000000000000000111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111100000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111110000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001011111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000100011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000010000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000010000011111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000001111111111111110000000000000000000001111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000001011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000010000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000001001111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000010001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000100011111111111111111000000000000000000000011111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111000000000000000000000000111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000001001111111111111111100000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000001111111111111111100000000000000000000100011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000001001111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111100000000000000000000001111111111111111000000000000000000000111111111111111100000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000001000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111000000000000000000000000011111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000010011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111100000000000000000000100011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000001000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000010000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000101111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000001011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000001111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000001111111111111110000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000001011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000001001111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111100000000000000000000100000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000001111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000111111111111111000000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000001000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000001000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000001000001111111111111111100000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010001111111111111111110000000000000000000010001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000001001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000001111111111111111110000000000000000000010001111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111100000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111110000000000000000000000001111111111111111000000000000000000000000011111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000011111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001011111111111111111000000000000000000001000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000010000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111110000000000000000000000111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000001111111111111111000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000100011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111110000000000000000000010011111111111111111000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000000111111111111111111000000000000000000001000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000010111111111111111111000000000000000000001000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000010001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000010001111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000001000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000100001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000010111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000011111111111111110000000000000000000000011111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000100011111111111111100000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111100000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111000000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111110000000000000000000000011111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111110000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111100000000000000000000011111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010000011111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111110000000000000000000010011111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000011111111111111111000000000000000000001000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000100001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000001000011111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000010000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000001001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000001011111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000010001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000001011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000100111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000001111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000001001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000101111111111111111000000000000000000000111111111111111000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000001111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000010111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000001000001111111111111110000000000000000000001111111111111111110000000000000000000010001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000100011111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000011111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000010111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000010000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000010000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000010000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000001001111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000010011111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111000000000000000000001000001111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111000000000000000000001000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000001000111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000000111111111111111000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000100000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000100001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111100000000000000000000100000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111110000000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111000000000000000000000111111111111100000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000101111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000010000111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111000000000000000000000000111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000001111111111111111100000000000000000000000001111111111110000000000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000001111111111111111100000000000000000000101111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000101111111111111111100000000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000001000001111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000001000011111111111111111100000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111100000000000000000000011111111111111110000000000000000000010000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000111111111111111100000000000000000000100111111111111111110000000000000000000010000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000010000111111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000101111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010001111111111111111110000000000000000000000000111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000010000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000100011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000010000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000010000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111000000000000000000000111111111111111100000000000000000000100111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000100001111111111111000000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000001001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000010000011111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000010001111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000100111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000100011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010001111111111111111100000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010000011111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111000000000000000000000001111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001000001111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000010001111111111111111100000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000100111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000001001111111111111111000000000000000000001000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000001001111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000001000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001000001111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000010011111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000101111111111111111100000000000000000000000011111111111111111100000000000000000000100111111111111111110000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001001111111111111111100000000000000000000100111111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111111000000000000000000001001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000001111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000010000011111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100111111111111111110000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111110000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111100000000000000000000001111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000010001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000011111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000001011111111111111100000000000000000000000001111111111111111100000000000000000000100111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000001000011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000010111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000001011111111111111111100000000000000000000000000111111111111111000000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111100000000000000000000011111111111111110000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000010000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111100000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000010011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001000111111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000011111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001001111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000001111111111111000000000000000000000111111111110000000000000000000001111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000001000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000010000011111111111111111000000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000000111111111111111110000000000000000000000111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000100011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000010000011111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000100001111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000100111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000001000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000010000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000001011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000101111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111100000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000001000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000001000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000100011111111111111111100000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000001011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000010001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000101111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000001111111111111100000000000000000000101111111111111111110000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000000111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000010111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000001111111111111111100000000000000000000100001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111100000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000010111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000101111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000";
	SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)		:= "000111100001010100111100001101101100101011101010101010011001111010110110000011011110001010000101110001110100100000010111101010000100001110011111101101011101111111101101000111110011010000001100001101101100010000010111100001001011101110010100100001101000011010111000010011011111011111010100010001001010111011111010100101011000101101001011110010001100101000010101010111011010111110000001110101101000110010010100111010010100101101000110011011101001100001110100110100111100101101100010111001110111110011101111101010011100110110111111110000010101101101110110100011111010111101101100100001101000111101100000110111011100001001011110100101001011101000010110110111101111100100101010110100111000101101000010100101001001101011100111011101010011001010110000111101111111111111111101110000010100110100100001000010100011111111111001001011001100110011001010001000010100010000110011111000001010110101101101111100000100100010010100100100101010100100110011000000001110101111011011111110011111101101001101110101000101100101101110101001101000100001110101111000111000101000101101000001111111101001011100111110001001110110110101101101000111000101110000011101010100110111010111101011110010001000111101000111011001101010001001100111000001011001111001110010101100101000101010111110101000110001100101101010111101100011010100011010000011010011101110111101101011111101101100110010000111111111100011110110011100100111000101010100000011111101011010011001110111111100101100001100100110111001000111011000110000110001101000011011000100011000101111011100100100010101010100101011100000110000011011100000011101001001011110001001000011110001111111110100000111101101011001111000001101100001011111110001010011011111111001010100111000110011100111001101100010001001100101101010111111100010001100100000110101100111001111001110110110111001001111110100100110010110101100000010011101001111100100101111101010010000111100011011100101001001110110010101111001000011010000011101111100111111110010001100000100011000001101111101000000100101011010010110101100001101001011111001100111011110110001001001111101101011100000100100001001110000001100110101010001010000101100100000101000110001000001011011110111101001101100100001000110100100010100011101010110100001010000001101010011011010011100111001100110001010011010100100100010000001011011001000111101000111111100000101011101001011110110100111100000111001010110000000011010101100110001101000111110010111101111100001001010011011000111111101001100101011100001011110001011011110011100001000011111010111000110000100101001100110100100111100101100100001100110101000011000010101000000110000110010110110110010000101100010101101101111111010111001101011101100010011001101101000011001001111101100010110111111111000101110001111110110011101010111101000010111111101010011100000010000100010001010000110110111101101110011101111110111100000001111111111000101111111001000001010001111010010111111110010000110100101010011111010011101100010101000101100111100011001010000111110101010111111110000001111110101011100010110110000110101011100101011101110111001011100011111011011011110001111101001010101011101101000111110111111000110100110000001011101000100110010111101100111011011001011101001000000000110111001110110111111000011001011001000100000100101010111111011010101101000111110001110100111010111010001111011011111110010100110111010110111011001110011010101111010011000001111110100111100000001100111111111100010001111001100110011010010010010011110011100101001011100101011011100000000001111101110001001100110111000110001011111101110101110010111100000011011100001001110111100110001001010001010001110011100101000001001100000100011000101100001111111100000000011001100011010100101101111011011101011110100100010111101000000011001100011001010111111101101111010110100101101111101000100100010101111111011010110011111110100111000101000110001010110101100111001110111010101011110001000100010010000100010001000001110110100100111111000001010101111011100100010110101010101011111001010010110001000010001100110100011100110101000011111010011111011110111010101111001010001111000000001101100110110110010110001000110010100100101011011111011000101111011110100111111100111011100111011110010111010001000011010001001111010000101001001111101111000111100111110110101000001110010011101111001100110101011001100110011011111110111100110111110100000100110000001010011010011000011101001000001100000110101001011100110111010000010101101100111110010010101110111100111110110001111111110010110001000110100001011101110000000000010011100010011100010101111101010110100111011010001111001111001010010001001111111000110111101011011111110101100000110111101100001010100000111001101101001010011100111101101011000001001001010001011000110010001101010101010100110110010101011110110111110010111000010001110111100001111011010011010010011011101011000110101110111111110010111011101010101110110001111100100000011100110011111001010001111011110001001101100000110000000101111101011011111110010011010000100010011011111111110111010000010110111011010000001100000101100010011000011110100010011001011100110101011001110110000000011110100111011011010100111101001001010010001000011101000000111111101000000110100000011000010000110101001001000000011011110011111011101000101100000111100111110000110010110101001110101011010001111110110000111111001100111000011101000110110000101000011011101001111100101101001010001010011100100111011011100101111011011010011100100011110101111111000100000001011101101010010000100001100011001010011111110110100101000000101001101011100010001011000111001100101101101010101010000110010110001111011100001000101010010010000010001111001111110001111110011011100011010010111001001101110100011101011110011100000011011000111101011000100110010001110001101100000010011011000010101111110111011110000001110000011100011110010101000110100000011000110100111101000001000101100100101000110000110100011001110011100110110100001011010111001001111110011000010001100100111100101111101110011111100000110101011110010101101111001111101110110011010010110101011011010010111001101100010110011000001001001110011110001100011101100011011000010000000111001001101100100110100100111110110000101010110010110101110110111001001110101101101111101000101000010001100101011000111000001000111111010010100111001101110001111011100001010010111010100010111000011001000011101111100111010000100111001111110011101010110100001101110011011101010011001111010011100000100010101001011110111101110001110110010111001111001000110001011001100110100111010000010001011111001011100100000110100101111100110001111011010110110010010010000001000010010010011111000100110100011101010111110111001101010100110100011011001101010101111000001111100010001100001000001100000100011111010111011011111100101111111100111101100001101101100111000101110100010001110010001000110111101000011000001010010111110010110101110010000100111011101001011110101111010101010000001101001110100000101001010101101110000110001100110011101100001110001001000100001100110011001101100001011000001001110110111010110001110010111101110001110101110101010001111100001101110010101010011101101000001010101111111101000001110101010010100100000000100100000010110011010110010110100000101101010001001001110000111110001010100001100010000001110111001110100010100001111101000111101100100000111101110011010000101001011111111001011010001110111000011011111010101110001101111100110010101001101100110000101100010111000111101111001000011010111001110110010110110110100111110001001011110110001011000011011110001100010101000101100001101011000100100100100010000100101101000110111011110001011111100101011110111011101010101010010010011000000001011100101010000110011101101001011000000001000111100001001000100011010111101000100101101011100001001001010001110010111101100011101100011111101110011101101111111010011111000101011010011000110110011010010111001110001100011000101001111100110000100100001011111001011000001110010110010011010001011010010000110010101011000110000111010100011011101001011000110001110010110100100100111111100101011010001111001001111011111001101000110100001110100100001111011011000010010101001111011010011000110110001111000000001111011010001111100101011110000010011000111111101010100110101010110110111010100100100010000111101100111001100001100011000001001101010101111111101000001110010100011010100100111110101001101011011110110100011011100111000000101011111101111011011110011011010101111010011101100010011100001110010101100001011010111101000110000111011000000100110011011111111011101000100111110011000110011100101000101001111100111101101000010110011101111011000000000001100000001011100001111111000100010011010001111101001001101111010010001010111100101101000100000110100011000110100011001001010100000101010111011100010110010011000100100001111001100111011010000110101010010111011001111010100011001101010010111110000111000110011101001101000011111111010100011001010110111110100011110101111000001011110111001101010100001000110011011110111010011010010101011110110110001011011011011010110001001101110010111011101011000010001110000100000011100010011010010011101011111100110011010010110010100101101000001010011100100001011100111010001110001101110101111010001001010110100101111001001001000111111110000011111101011011011100010000101110110111011010010000111111111111010011000110100010010110010110110100011011111101000101000110100110100111001111011100110001011011011100111110101101000111101000001000010101000110000000101001101011010010111010101011011110001100011010001010110010011101011111011010110110110000100010010110100101011000011101111011111100111100011010010001100100010001101011111010111011110111000000111110011010110011101011110000000010101010000111111000000101101010000111011100100001101010011100111011110010000100010111011010001000000010101100011001010001011100111100111000000010011001101011101001110111011100111111101001011100101100110001111101111111011000011000101101111101100111110011110000101111100111101011100100011010011101110111000101110010010111100011110101010100111001001110110000100000111100111101001010111011011010010001101111101100011010110011011101001110111100100011101011110011100011111111111011000000000110110100000001010011010101001011010110111101100111100101000111001010100000010101011110011100111100100101110011001000100001101110100000001110101001000000100101000000101100000111000111111110111111110001011110011010110001001011110001000010011010000111101011000110011000001101111100000110011110010010000011100111001110001100000110000110111110011011010111010111001110101100011001110010001100011110000111100111110100101011101101011100011011011111010011011011101101000010011101101111110110011101111111101010111101111110101111110000011000111000111110000100001000111010100010111110100111000110011001101111101011010000010111111011001001011000011001111000101110101111110001010001110000101001001110110111100001111000000000100111100010111111100100100111010010110000010000000010101011001100010011010101100001111010010001110011011001111001011001001100010100101001110011101010101111000000010011011010100110110001000110111110100100110011000011100100010110011011001000001111000111010100110011101110010010101101011000111011001100011000101001100110101111010101001111100111001100000111101001001101001101001010110010000000110101010100101000111110001001001010110110100110000111001101011011001100110110010111111110001110011111001100011001010100010100110010000001000111001110000011100100110101010101110111011000010110110101111111011111100011100010101110001010110011011011110010111001110101100100110111111010001110101010100110000001000000110101000011010110100101111000111111101100001000111010001110000011001100101100001101100100011111011100011011110000000111111110001010111011110011101011000110110101010001011111010101000010101011111011110010110101001010111001001001000101011111000000011110100011111001111011100111100010101000110101001001100000111010110110110111011001101011011010010010001110001011101100101001110101010100001101000000010101000101000010100011100000011101101011110011100000101110010100110001000111101011101111101110001010100100110111111111001010011101001000110010101011100111001100100001000111111001011100000100001010101000010100001100011100100100000100001100011101010111011110010111110111011100111000000000111000011101001001100010101100111101010011000011000001001011011111110101001001100110110011101110100111011110110100101100001000110001000000110001000111011000100010011111010110001011010000100000010011100111000001100011111101010010001011101110110101000000001101111000101010110010000001101101100111110111000101100011100111001011000001010001010111101100010010000010001001011101111011001101011000010110000110011001011000111011111110010000001111110111110000011100101011010011010101111100011111111011111111011111011000110010010010011111001001010111110100011111000101101100000001011111110111101100111111010001110000100110011011011110001101001000010111111100101101000101110000010010110000110110111000111110000101001001010000001111111010111101100100001100110111101101100001111110111100011001101110100001001101011110100101011101001000010100111111011100100101100010000110100101011101010101111100101101111100000111011011001011101010100101101111001000010101010111111011001000100001110011111100111001001101001010110011100000111010011011011100111010010010100110011010111001011110101010000110001110000010101100001011101110010010101001101110101100000110110011111101100010010000011000110110010010010001101001101001010000101011110100010000000010011001110010010100111010101100101000111101110000010001010010101100101000011011010100111011111010101110100110000011110101001011011010011110001010010010111011001110011111010011110101110010011111001011000101001001110100111011110111110011100101010000011001100001001000001000001001010010000101101011010111100110010010100100101111101010001111101001100000101100011101101100101101101010001010100100110000100010010000001101100010001101000001010000010111101011111101101011100110011110011101010000011101101101110110011010100010000101111001101110000010101011001111110110000000111110010000101011011111111111100000011001101010000010011001111011110001001010111000110100111011000011011100011011001110111111101011010111000001101001111110110011100111110101100011110111101011010011101001100110101101101011010001101011100000100101000001100101011010001011101100001011110000011100100100001001010001101110101001110101111001000110001000001111110101000010001101110111110000000011011011110000110000101101001011100000011111001011011001101000100001110110100000110000011111101100100101100000111001100110010101110010010011001111110010010110111101110100111110001110001011100100111111001111010100001110101011010110011101110111100101011011001111000001101010101101001010001010100100010100110100110010001111101110101010001000011100001000001011110000111001000000001011101100111111010101101110111011110011011100100010110010011000100111100011001100011101011000000100011101110110100001101000111010101100100010110011110000010100111000110110110110110110111001111001000111100110000011100101101000100110110100010000000010110111101011001100010001001000100011000000010101101001111010000100011000100011111111111010000000001100101111010001101010010110011010001001011101110001110111110100010011110010001010101001111111111000111101110111001010111011111110000000001001001101100000101101100000011100111111000111011001010110100111110001100101000010001110011111001010001110111100001100010110100001000100000010001111011000010110001001000100000110100110101110010100010111000101011111111101010100011010010100101011110010010101010010110011011100111010101000101110101110101101101011111010011000110011011101100010111101011101101001110110011110111010010000100100001011001010101101000001111010111001001111111011001011101111011011111010101011100011111011000111101110110001100011011000101100100000110100001100010111001100000010011010011011001111101001101100010001000110111110011010101010010101001101000101100000111100011000000000000101110100001101101100001001110111101010110010100011111000010110011110110001101010100101111011010000011110100111001101100101011010010011100111100100110111101001011110101010010100110110011111100010100100100100101100000111101010011010000011011111100010101110001111101001001111110100010110110111100111010110001011100111100101001110010000010011111111111000000110101001010101001011010100011111100011010011010010100001100110001001000011111000110110011111111100101111001011011010100100011100000001011010110000110111100110011111110110110100010100011001111001010100011111000001111100101100111001010100001000000000010110000100100111000010110011100011001110110100100111110010001010000011001111010110011010010011101000101110000111010001000011001110000011011111111100011110101110110110111100110110000010111011010011100111111111000111000010100101011000110110100110010100000111001001011000010000001000100100110011101110100101111011100000101110111011111011010111010011111001001000101111010110000110110010110000110110110000010010111110001001001111010011111011011101001010100111100001000100101001110111001000101110101000111101101011010111110010101101100000011001101100100111110111100110110100111011001101010101100101000011110111110101110011100111110110001101001001000011010111001100011010000000001001001001110001001111010001010111000111110000010101101110010010111010001001000010101111010100011101110000110110100111000111010100000100110100110110101000000011110001000001100011100111001011101110001010001011000101101000000101100010000100101011000010011110001000001100011111011101001000101000000011010100111010110010101111110001101101000100001000010011101110111111110010101101010100000001101011100101101010000110000011101111111110001111101000100011111100011101101100001100010101101010101101010101100101101100101011101011011101101111000010001011111100000001010100010011001001101011011101010110101011110101111011010100011011001100110101111010111110000010011011101000010011110010010001000111111111010101111010100111010101100010011000011011101100110011100110110000000000110111100010010000000110111000100101001110100011010100010110011101110101101101010101101010101100000011101111110001100000100001001100011011010010111111101100110000011001011101010001000000010111010010111111000000000001101010000010011101111100100111000000101010011100011100110001001011111100100011000111011110101001001000111110011000110111100010001001001111001110100011000101111001000011111001010011101010000101101111000001100011101111001011001111011001101101001110011111101101000001011011000111001010000101100111111111001001100010000000011000101011100000111010010100110100101111101011111001111000101011100100100101001000000011000111111110010101110001000110101100100111111011111000111111110010011010110101011000001110101011011001000000000000000100000011110110010100110110001001010111010110111110011001010110110011000101000111000000111010000010101100011101111000011110001101011010011010010110010011110111111001000011000010110000100001011011110010110010001111001011010110000010101100110101011100110011100011101001101001101100011010001011010010010100001101010000011111111111000100010101101111100011010111101010111101100001000011010110011010001001001000011101111111011110010010101001110001000110000011001101011011011010000011111111111000001100100101001010101110100011001001110000100111100101111110011110111110100110101011101011011001011001101111111110001101111111011011010011111100100011001000010111100111100011001001010000111111010111101101111011010011011111000111000010111101010110010001100100001110010010111111100001011110000001010110010100000010110101101111101101011100101000000010101101011101110011010110001100000011111001100111111010111101011111111100111111010010110111100101101010011101110100000001111101001111011111011001010101010111011001111111001010001000101011010001010001110011010110000100100100101100111101100101000111000011110110001100101010111011001001101010010110000110111011001111111001000011100100101010000011110101100000001100111110001101001100001011110011010100100100101011101000101000100111101011110011111101011101110010100110111101110000110111011000111111100100101110100001110001110101010101101101111101010010011010111000000001100110010110100010110110101110000110000111101100001011110001001001101000011001101110101010011100001110001110011001111000011001000101001001010000100000100001111110010010110011100111100111011111111001100010110001010110100111100010011001011100000001101110010011000100001000010011101110110010011011111011101001001000011111111101101111011001101101110100010011010111000011111000111111000000101001000101110010000011000100011000001111011110101000010101011100100000000100101111011100110000100101110110110011111100111010010010100011000011011101100111111111111100001010101001110010100101001101000111101011010010111000010110110101011010001100000111010000001011110000010111010001111111110010101000101000011110000100001111100101101101001110101010101110011011101010110111011101100010100001001001111111001110000110010011011100111101101010111001001101110000010010000100010001111100110111001101111010110110100011100101011010111101101110000001100011011110101001011010101011101001111111011111010001110001100001101110111111000101110000101100101000010100011111101011101111000111111101111111110100110001011010101010110110111110001101010011010110100110001101100000011111000010011010100100111101100001010110100110110001100100011110110011101101011111100000000100001111101010010010001111010010010001010000001111001011111100111110101010001011010100111110010110011000001110111100101011000010011100111101000111110010000111110010110110011100000111110101101111001100110100100111000110000000111100010001110110111000000100111011010101011100111101000000101100110110111011101010010110000001100110100001000011011111101001000111101001001011100000110010100001011100000011111110010010001101011011011010010011010110110101111010001011110100001110111001100101100011001100001010001000010001000110111011111011111001001010111000010011111001100000110010011100110001101111001110010101000001111011100011100111100100011011010110100101010010000010001011111111110001100001011001011101001011111011110110101011011000011001011010001001110001110101110101111011000101100010100000111001111011000001000000010001101010010011001010001001111110000001001001111110000011110111101111101001110001100001101000101100111100111000000110010101111111010110100101111110101111101010111000100001101101011110110100001010110111111100101100101001100111001111000010010011111100010111111011101010011111001011001101000010001001011010010011101111001001110000000001000100110110111011101110101010101111000000000000000011111100001000100001110110111000110101011110100000001001011100110000000111111111001010110111101110010001001010001100101111001010000100010001000100011110001011000011101000010101111011110111100000101001001011000110100111011000010001011100110010101101000101001001000011000110010000101010111010001101101101101110101110011100001000110011011011010011101100000010100011010011010111100110101011011100100101101101111100101010000000110001010001011011000011011110011010101100100010001111010100101010110100101011001100101110100100011101001010000000100101110111001100101100010001111001001111100011001010011011011110011101000100111011001011010000010111000011011000101010111110010101111110110100001101001101111111110010010101101111100100110101000001111100110011100100001001011110110110000000011011110101001010110110101111010000101011111110001111111111001110011101100111010100001111110110100000110001101001100010001001010100110010100000100010010111100000011010111100111010101010111100111101000110000001111111010001010100011011001001111111101001100110011001101001011010010110001110100010010010100010110001000100110000111011110101100111101100011011110111011011101100010010011111001111101111011100100110000111000101000101101110110101001110111011011001010101000000001000101010011100111110010110011111000100110111010001000110100100010011100001110111100110001011110100011001111100111010100100110010000101101111100111100100100101011110001100110010001111010110010101001000001001000101010111110111000110011110110100110111011011110101010100000111001101000101101100001111011001000000011110111101110111001100111111101110010111001100011000011011110100110011011100010010111101011101010101001011010111111100101001011111110110111111001011011011011011110010010011010011101011000111001011111000101110110011001000001111111101101000000100000010011100010001110110011011101000101100101111011111100001000110001100101101011110111010010101100011101011101111000010010001011000000000101100101110000010000001010010110100110110111001100001010010010011111101001101011001001110110000011101110010110000011101001100000111001000000111110010011111000001111111100001111101101010001101011000101110110110101001010010001010010100111010110100011111010110011111100101001001110011000001101000110101000111101110100010100100100101000111000010101101111101010010000111101100010011110001001010101001010101010000101011101100011110101010111101111000110011111110100001100101011100110010000110010001000101010111100101001111011101011111100101000110001001010000010000111011000000010101000000000100100010111000100010000001011010110000110101110110001111011001001111001000101011100111101000001100010010101110110011111110101111010000011101011101001010111100000011111000101111110010001000011101110001111111000111101001100001111111111101111011100001110110001011011000000010100101010111101001000100100001110000101101111110100001110000011101000101100110000010111000100111101011000010001001110010000101000000101010110011010111010111011000011110001100011100101011100000000110011100010100000111100001110101101010111101111101100001111010000000110110111011101010101101001100100101110101101101101010101110110100010110000001001000111110011101111101100001011110100000111100101010010101001000000001011000001010011010101011001111111000100000101101111111000111100101001111011110110101101101111011000011010000101100001011010010001100111111011000001011100101011001111101110000000010000110000000110101101101000010011111101100010100110011011101001011111100010011100101111101110110001101101111101111010110000111100001100111101011111010010111110100101111011001111100110000101100001101001001101011010101000101001010001100011101011100110100110110011110011001110011000001111010011010001011111000000010010011111011010111100101011011111000011110101001100111100111101101000101000001111011101000100101000000110000100011010000000001010010101100011100101110001101100010010111100011100100011000100001010001010110100001101101110100101110100010001001000000011001101100011100110000010001000010101000100111110010101100110001111100111011100100101110100110110100110111001111000010101011010001011111110110001100100001000111100011011000110110011100010010100011001000001100100101100001000111000101001011011010111011000100111110110000001101010101010000000010110100110010110101010100000011000000000100110001000011010110111111000101110000100110111111011111011101110010101000110000110001110101100110011011110110100100100000111100011000111001110110011001011010010011001100001100100001101100110000001111011001011001110101110010101000010101011011110111010111101100001100011010001111001110100000000001111011010110111111010011010010011001001011011010000100101101111011010100101000111111110011011001010110110010001110111110101101111111010100100000110010110110011001001011011001011001011100100100111101011111000110100001001000010111111111000111011010110011100110010011000011101010111110010000001111011000010111000011000111000001100000111111110101010110001100001001111100101001101010000100011001011100001011110011001111001101011101011000011010011011100111101001001101110101010111010101000011110111010001010101111111011111111010111000010000011111101110100101110010001101100101010110101110011110111001011011110001110001010001111011010011110001110101101111100011001001110101111000111010100110001111001101100001001000000010011101011011110101111101101010110010100111001011111111000001111001111111010001111101100101111101001010110100101011011011011001011000101111011110010011110000011000011011000000011111000000111101100001100111101101001111101101100100101111010101011001011001001000010001110101100011011001110110000010011000000110010111100011001000110111110000101011101000011111101000110000000110011111011001110110001111011011101110101110010111110111100000100011000011011101001110110011101111000100110111001011001011010111101010000000100000010111001111001001101111010101110111010111100101110000110101111101100000100011111001000100111010010000010001001011101010100100011001000101011010100110000101110010010001001001111001010110010101100101010101111010110001010000011101010100101110110010010100011101001100101011111100101000000101111011010001000000011110111110000111111000100101100110010011100011001111111000110101011101000101001111110111010100100000101100011110101100011111100101110010001010010111010011101000100100000001100001100011011000011111100101010111111011111111010011011011000010000001101001010101110010010000001111110011001111100100001001000010101101000010010010101000011000111101111000100110000100010101110101000000111010000010111000101111011010100100101110111100111100000100110010000011011001101001111110011011101111100101000110001101010011111110101010101101101100010010100000010000011010011001100011110000101101010100010111111111000001011100100010011100001001111101011001000000111100010000101001111001011011001101000011111100100100010000001011101011000011111000100011000001010101000100011101000000111010100101000111010111010001001100010011010100000000111100101000000011101110001000000101001011111000000001101111110111000001110011100011101000000100110101110010111101001001011100110100101011101101110001100110001001010010101110111011011101110110100000011100100111010001011011001011011011110111001110101100111001011111010011111110001110111011010000000000101111100100000001011010101111010011101011101110100110000100111010101111100011001011000111100111011001001111000000010000111101110110111000001010110000000010110111111110011011110011110011100011100001110110001101010110010100011010110001011011111110000111101011001000111000110011101100001100001010010100001000100111011011100111001110000001010001100001100011011101100001111101010010001010011101000000111110100010001001001100100001110110111110101101110110100001010100101000111100100111011101111000010001011110001101011011111101101101101101011000011000111011010100101010101101000111111001001011100000110001011101001110100000010000101010001010101110010001100110011010111110000000110001011000001000100011000101111101110111011110010011000001110101011111101101100100101110110010000111010111111110000010110000100111000000100100001101010101010001111101100000011101010010001101001010100101011110101001111100110010010111011001100011111010010000110110010011000100000101010110110011011010110011110101101001111111001101100110001100100011100000001010011111101101011000100111101001011111100101101101110110010000100011110101011111000101110110110001011110111000000001000000000101011011111010110100011101010110100011000100110101111100111000000101000100111111101111000110110101010001010001100111000100100000010011001000100110011001100010011000010100011110011000001111011110110010000010011110111010110011011100100001100111100101001000100101110111100110100111101010110000011001010100101110111001001101000100101000101111111111001101110100000011101111001110000111111001001110011010110010111001001001010001101111001011100111100100001011000011110110001011010111010100010101111110101001110011001011100111001000010101011000010000110101111101000110001100000110010100000110010100000010011000010010111001111000110111110101110000010010100101001010011100111110010001001110000001110000001001111010101101101000110001011011101101100000011110100101011010101101101010010001100000001110100001001010111010000100010000100100000001011111111101101010001110011101100100010000011001010010000001011011101101010110110001110010110110000100111011110111010111100010100110101010011010100110000000111010001100111110010111111100011011100001101100101011111001001100101011011001110001011011101101010011011011111110011011110011100011111011111001100100111001110111011011010011000101010110010100000100111111001111111111100000100011011010110101000100011110011010101101110010010001110001110100101001001100100000011010110000110110110111000011110111101011110001010010010110100101111010000011001101001000111000110011001010011010111001000100111011011111011110000000111100000111001011000001010010010101100011101011111000010001100001111000101111100010101101111000100001111000110010000010101001010110001100011011001011010100001011010110101010001001001010010110011001000100011101001011111000100111110010000110110000011011001011100011011111111111010110011110110100001111110001001011000100011110111011001011000110011111001000101001011110101111000001001001011111110010001011101011110010000110101001101111101101110110100101100000110000011111101101110010100110011010100010011101100110101001100000100010100101000001111010011000110101111010110011111101001101100000001000100101010010100000101111010110001101010000000111100001101100100111001101010000011100100000011100000001100111010110001000101000010101111010001011011010010000000101000110111110110011000100101100100111101101101101001110011100111111001111111101111000000101010010010001110000010010011011010010110110001010110100110110100100100100000011101101011101011101100011100101101110110001101011011010101001001111111011000100111101001001001100000011001100110101010101101111111100001110001011001000110101100110100100000010001100000011100000001111000101110111100110110100110100101100110011101000010001111100000111000000001000011011100010001111011110011110100101001110100110101110010011110111111000000110111111000110111000000110000101100100011101101011000000110000010100010001101011100101100010010110011011101001010100100011100101110010111010011101100011100000001011101111001100000011001101111010111111001100000010100101101000111111110110110111101110010001011011110110000100011001100000101110100011100011000100100010111110110110111100000000111101011101101110011000110011110010011011010101101100111001011001011001101101010110011000110010110111011111011110011011111001001111010100011101111110011100101010111000100101001001010101101100010011100010001110010011100010100111101110111011100001110111111001000010111100111110011111101011011011111011111011000010000101001111010101001101101101111111000111111011010011010101111100110101010010101111000111110001001011010001111110101110110111110100110001011000100001100011111110010011011111111001110100111101010111110010101101101010101001111001001001101101110011011001000001100000000011101001110100001011001101111110100111000110100011110010001001001001101000010010000011110011110111011110010111010010001001110101101111111011110000001100011111011000011000001110001111000101010010010110010000100000100011100100111110101011011011010110101110100000101011101010001010011001010010000100111001111101000001110011110000101111001110111101011000101100111100001000000000010000111011100011101001011110010101100101100011101111111110100011001001101001111111100011111101001111000101101000101111101000110111110100110011110110000100001101010011101101110100100111110100101010011101011100000100011100001001010000111010001011100001001010000000101110001110011000101011001010110101011110110011001010001011011000000010010000010111111111111111111100111001001001001110110000001000001000110100011111111011100111010101000111111010010010101111001100101000111011110100110110010000001100010110011100100010100111010000111000100101110111111011000010100001010011101001110010000010000111001001110010111101010011110111100011100110001100101000111110010010000110010000100000110011111101011000110100100100100100110101101011110111000111101011010110100110010100111100111111011010001001100111110111101110011111100100101100000111100001011110010100011001110110100100000011001111001101101010000010000000011110000000100011110010101011001110011110100010011000100010011101001000100111011011000101110110110101100110110100000101100100001100011100001000000111110000110100000100000111111110110011101100101101110100110110101110001101100110101111100000101110110100001011011110101101001010011101111011101110001000000100101000011011111100110111011010010110000101010010011101101010101110010001101100110010010111101111001110110101100100110111100000011011101111111011011011111000110101010101000101110111000111110000100100100100011011100010100110111110011100110100111010001011001110001100010011100001101001100110100000010001000101111011011110000100000011000001001011111001111011000111000000110010011011010001010000001100111100001000111110001110110101100010100100011011111110000100011110110001011001110101010000001001011000010010001111100010101111000010001010100101111110001000000111000101100011110111100100110111111011100001101101101011101101110101010000010011001111001010100100011110111011101001101111111010100001110001000101110111110000110011011011010101111101110001001110110110110011000100011101111110011101100111010110111111010100110110110001001101101011110000010011110000110110110111000001101000101011010011011000110100010011010101101101100111110100001011101100000100101111010100000010110111111110100101000110001011100101010111010001101011101001100111001110000100111101100111101110110010101011011000110111110000010101110000110011111111100100000110010001010011111010110000101101001100000100011100011011110101000100001010010110101100011011101011101010110000010010011000001010010011000010100000101100110100001110111001100000111011101000010101000101011100101010011101010110111101101010010010001110010000000100111011010011000101011001111011111111101101011110001010111010101011001101010001001101001110011111011100101010101111101110110100111011110111111010001111010000100001110011011001010010110101110110100101011110000001101101011001111100111001000111100000001000010011101001011101111001110111001110011101010000001111100100101110001000111010101100101111000011010010010101011101001111110010100101110101110111001011001100011110011000101110010000111110101011010011110101010101100110101010001001110000010100010000000010100101101111110011000101101101100110111000100101101110100111101000100101010100110111011000010000010100111001111110001100001101000010011010101011101110110000000001100110011101010011100111010110011000100111100111001010110011111101010100011011001000001001010010000100011011010001100001111010100100101000001100110100110010111001001011010000011011100111010011000110111010111100111000000111011110111001101110001111010010110011000000010011100011000111110110110000101001011110100011001110110011100011101111101000001100000111011011100111000001011111011000111110011100100011010000010110010000100011110110110000011110010010111111011100110000000101011101001111010000100101010101010100111110011011101010010110011011010000011001000010100100110100000111010011001110010100100111110001100001000001110110001100101101011100101110010101110101101011111011111101001101000110011101001101111100001011100001100111101101111010100110110001101001111000111010100100001001110110010010010010010100000111111101000010010010110011110011101100011101000111100011010010000010100111101010000111011101001011101100100000101011100001000100010011110011111010000100111000110010000110111011000100000001001010001111000011011010100011110101011100111111000010100010110100110000110000100001000110110110110000100001001010000000110000000111001011110000100110101000011010110010111011101111000101110110101110100111000110101011101011011101001101000011101110010000001011011001011100100101110000011101011010110011111001001111010101110100010101001101010011110011110010100111110110011100110111010000000110100101110110110100110011000100001110010001010011001010011010010000110000001010000000100101000010001011111101110110101010111100110101011001101011101001110101011101001010110110001011100111011101100001110101110100110010000010111111100000011000110000110101010001101101110111010101101101011110011110101110111111010001110110010100100011111001111001111111010100101011001101001011011111100001010100001100001000101110111000001110101111011011000000001110010011011000110110001111101111110111001101000110011110000111100011100010101110010000100001100111100101101110001100001111011101110101011111010101000000111001100001011011101100110011010000010001100111000111111101111010000010011000010011011100101101010010100101100110110100110111110110011000000110001001100010110111001110011111110000010100000010010001101011111110011111011011000111101110001001000001010110001110010101100010011000110110111011110011100111011111001111111000011111000101100100101100001100100001100100100110111010010001110000001001100011110110011111101010101010100001000010100011001111001001110011000011110001011101001110000111110110101101111001010111010110010000000001000010100000111101001111001001000110001111001101101010010011100010110000001111000111101010100111111100001101101100111001101110101010011000111100000011010011000000011000000000001001110010011001111000111011100100101001110110101111000110110011100001111010111011010111011010000010010100000011101101000110111001010100110001101000110000000110101110100111101110011010000110111000011001101110011010001110111100000010110111011100101111001100110001111110100100001000111010101000000100101100001101111111101101110000010110010111000110100100010011000000110110010000100111001101100001101010100011111111111010001101000111101001001101010000011101010011111101100100001011000110110001100100110111101101111010011110111010011101100100111011100111000110100101000000011001011101000010100001010101011111101001110111100100010001101110100001101100000110011000010101110001010001110011000111100101011010001110001110001111001110110110010110101111011010101001001111110111010001100010010010000110101110011011111001000000111100110101011110110011000011111011000101001011000010111010111010100001001110101001101100110000000100001011111000101001001010000100101101010011101011110110100100010111011000110001001111000110100110100101111000010101010001000010111000011001000010111010011001101101110101111011110110101000100100111101110101111101010110000110001100011101011100011001101011000111110011011100111010000110111100010001011100000100101000001110011011011011001001010100110010100000011011011111001000100000100011101010110011100000001010100101000010111101100001011010011100011110111010010011000011111001111010101101100110110001101001111110111011010000001000110101101110100101110010101100011001011111000111110001001011101100101111100011000110001011000001011101111001001010110010000110000111011100001110011000010111101001101010111110000010000101100000100111100111101111011110101000000011001010011111011000111010011100101001001001111111000010100010100011101001001100111010111000000010110110001010011111100100000100010011101100100110010011011111000011101100110011011010000101111001001110111001001000110001110010001110101011110111100001110101010001000100011001110010111111110111000110101110100101111111101001001101110000010011101101110010010111101111011111001110011111011111011100101110011011111001010010001100011100001001110011011011100011010111101000100000111000011010100100111110110101010111110110010111001100010100100011111011100111101001000010111101010010011011010011101001001001001111101110001010001001000111111000011011000000100100000100101000101011100001101110110001000010001011101000001001010011100001000111010100010001101000010010100011011111001000111110111101111011000110100000101100010011110011001101010111000111010110010101011011010010110000010101100100101001001011011010100111000011101100001100000100001000100000101110010000010010001101111011000101101101000110111000100010001110110010110100111001010110000011011010010110010001010001010011000100011111000101111011010111000010010000111110101101100111100111101010100111100011110111011111010100100011001110110111001001000110100011010010010101110111000111000100101100110110011011001100110001101111001011101001010101110111010000011011101000011111111110011101010110100010100111001110100111111010100001110110011010011010000010001101011111001000010100010000100100010000001010101011110000111011011110110111010101100111101010001110101001110110101010001110011111111000000110011101010101000000011000110110010010010111111011010011000001110100011000011001011110001101100101100010101001110111110111110111001111010011011100110100111111010110100100101011111000001110100111110010110001111101011100111010010011100111001010001110110110111001011000001010111000110111011000111100010000110011110110101111111111001100100100000110111011110111011011011111100110000110000001011010011010001011011101110100100101101100100011000111100010001011010101101110111011010101010000010100100101000001101111010100110011100110010101000111101001000101011011101100001110110110111011010011000111010100010110110000111001001101101110101100100101111010111001111110000100110000001101100111011010100011001101011111000001110010010001100010011110101101100010100100000111001011011000001100011111000001111010010101001011101001101110101100101000100000001010110010100111011001101000011100011000110101010101110101010111111011000011010100110010001100100100111111011111101100110111101100010110010110000101100101011111000011101101000000101010110011110101010000010000011111100010100111110001111011000100001100010011110110011011100100010010100110100100100100100101011110101010011011010000000111011000011000100110110011010010110101000100010110000011111100000010110101110110010010000000010110100011011111001100011011001110110101001110000011100110101010010100001001111011010110111110111001100011110101010110101101111100010000110011011111100111000000010011111010100101100011000001101110100001001101000111100000111111001001000010110010011001110001011111010011100111101111011001011011111001000011111011010001010011101110111110010100000100010010001111110010001010110011001110100001110100011111011100100111111110000101011110011000100010110101001110110111011111111000001110000010010110000000111000011100100011000101100101100010110101010111011101100101101000011000011001101101000001010011000011111110000010100011111001011010101010010001100101110000010000011000110100010110110100011101010000111011111110010110001110101000101011110001101001100011100101000010000000011001100110100011100001001010100011111110011001000010100110101111111001111010101000101010110111011010001101010011010010110101111110101001011111110101010000000111100111000011101110111011000001011100010110010011001110000111110110001100111000110110101001001010010010000110110010011000011011110001011010111111101110000111011010101010101011000100001100111011001110101111011010010010000011001111011011100110001110000100001101010000111011001101001111111000100011011111100001010001111100011011110111101010100111111011101011111110101000010101011001000010010110110101001111101000011110111000000111101100000111001100111011011000100010010100010010101111011101110000110111001111111101001000111100000011101101100110011101011010100001000111100011100110110111101111110101001000101001101111101100101011110110111000111111001110001101010100000010101011010010011011010101011100010101011111011111011011000101000011011010001010110110011000011111101100000110100111100001111101000001111010011100111011111111110010101111111001000010100101000110101010100111010111001001101100000111111010010011101110110010010001000010100001000100100001001101111110000101101000101100111100110010001111011000011110001011000001010010111101010011000000000101110100110000110110011011000000010001111000100000011011000011110001001100110011100011011010111010010111110011100001111100111101011011000010001101011010010101000001101111100110001110111100111010001100011111011101111000011111000101110111011001100100100101001001000111111001011001000000110001110010000011101110100001010001100001011111011001101001010011101001100011100000001000001101010100001101101010011101100010010011101101110011111110101010100001110001111101101100010110110011111100101111100110111101011100100111000101111110011100000100111101001111100000101100010011010011110010110111101101000110010001100111011100110010111001001110101100010010111000010000011100011011010011110100111010001100001100101010001100011101000001110110001010001010001011101001011100101011011000010011100001010011001100111001000111101000110110101110001110111110001111010011010111100110110000101111010111010110011000101010100101100100001000111101100001001111100100100100010101110110011111001001001100001110100100111100111011001111000111101111010110010100001001001110000101010100101101010100100111100100100010100101101000110111010100010101100110010110010101010101100101011011000010110011000111010101101001111111001110011010010101011101001100111010111000100011001010010101001010011000100110011011100101101111101000000101110101101000010100001101111001001010110000101011001000110000101100111010001000011001010111001011010110111000110111101110111010001111100101101010101000101011011011010110000100100100011101110110010110001111001110011000010010101000001000110010100100010110101001011001111000111101011010111011000001000110101001010010010000100110101110101000111001010000100101010111000011011110000111000111111110000110101110010011111011101001110010100001101000110010000010100111110100100111111111011000100101000011111100010011111110011000101001011111000111101111101111001100100000101101111001001100101101001000010111011111110000110110010011011101111001110010000101101110100000110100101011001011110110011001110010010100000001111001011101111101011100110111010101001001100011001001011100100011110010001010101000100001111101100100110100010011010101001100110010011001110010001110110000010001011111111001110000010000010101000000011111101011100111100001011000001000001000000010101110111110000001100101110110100010011000001101100101111111001100100001001011101110001101101111001010011100111010110110100100001111010110100100111100001000011100100101000111011111101001110110000011101100101110000111001100100001110111011110101001110011111100100000011000110011010011011110010000100011001111111101001100001101111000000010101001111111010101010100101000100111101101000011010110111101110000111101000001101101001110010100011110101011100001110011100111000100110011110010110101100010001011010011001101110001111110000110101001110010110000001111101101110001010110001000110100010101100100101110011001111010001100111111010011111100111011100110100110110010110011010100100110010111111111001010100110011111001110001101011101100110000100111111011111111001110110010101101001111000111101011011001000001110000111100010101111111000100010100100110011101001001011011000110111101001001110001001110001010001011111100001010100110000110001000110100100111110100001011100111101111001101101100101000011010110100001010100011001110111110101011010001101010101111110001010010000101101000110010011011100111010000011100101011111011110111000010110011100100100100000111001101100101100011101000101000111100111110101111010000001100111010100100110100100011011110001001110110001000101111101010101110110001101110011000100001101100101101000101111100010110101110001001010111100001010010111100000100111101111000101000111111111000111001010010111101001110010010110000110001010101000110011100110101000101101010110101010101001000110101010111010101100110101000111101001111111001000101110100100011001100111011010110101000110000101101101000101101000000000011011101111110011010111000110011100011111111000001100011100101001101000111010010000110100000000101100101010110101101100011010110010110010010001001000011110011011110100110010110110101011011010100011000110101010011000010001111001010100011000101010111110010111011000100100100000001000111010100101111110111100111110111100010100110110101000100001011100101101010101001101000111100011100010101010110001100101001111110000100101010110111010011001110111100001110101100000001111111111000111111110100100100011010010101001010010111011100010000101010110111010001100101011000000111011010000011000101110111001001011100111101001000100001001011100000110101001001011001110101101110100011110111110100101100010100001001111000010010011101000110100011000100100001111010011000010101011101011100101111010001000011111011101001010100100000001010000100101010110001110110000000101011011001110011100110101011011010001100100000100011110000100111010010011111000100001000111000110010101011111011100011001001111011110110001100011111101010110011110010000101101011000010101101100001110011110011101011110100010011110101110101010101001110011110000111110011111111111010001000001001011101000110101101100111001111100001111111111000000100110001110010010101111100110001010101010110110010000010011110110110001100010011111110011011011011001111001111111001111110100110100101100100001001010011010010011001100101110000100001010000100001100100111001010100110010011010110101000000110000001010011101011100001111111011101000000001100110010011110111110000100011010100010110111001110010011110100101000100101001100101000010101101111101010100011010000010110111001001011010100001001001101101001111101000100011101000111010110111101001001001000101011101011101001000101110010110001101000000010000010011010101111011011100110011010011110111001111001001101101011110111000101110011001101001011100000011011011010100001000011000001000100000010000001111100000010010101010000011010111111111111110000100001000101010111001001111111000110010001100011000011110110111000111110000100101010010100011100110011101010000010010100011101001100000000001101110010110010110011101100100010101111001101000011100001110101000110000010010010100100011111010100111011010011001101000000000011011111101101111000101001011111001011100101110011101001101010001101010110010010111001010010010111000100111000101000101100000101011010000001011100011001101100110111111000101010110010100000001111110101100110111101111100011000110000100111001111111001110101000011101110111101010010000110110000111000100110100110110100111100001110010100010110010011000000101001000010110101100000001101100101011110010000110011011110111000010111001101101010001100101110001000111010100100100100001010111011010111001101110101100101010100011011111100011011000000101110001110100111011001111001110111011111010100110011011110111001000011110111000100101110111001010110001101010100100101010100101000000101011000110111011000000111010100110000101011001110100001011010111011010010101011001001000000001100001110101010111011111110001010001110000011101110101111111110100110111000101100001010000000110111011001111110111001110110001011000111111001110110000111110100111010110101000101010110010011000111011111101001111011011101011001111101110111010111100100001010100101111001100110111010011101101010111100010111111011110110000110111001000011010011001101110110011111111011001001010100011011100001110011110101101010111000110100000110101111010011001111110110111111000011010101000000000111010101100001101101010101100100000111100001001010111101101000111010111011010011110110000100001110011001111011101011000111010110101111001010101010010101101100100000111001110111100010111111011001010100100101001010010101110001000000001001010011101100110100000011101001010101110011011110101000111011000100011000100110011100000011100000010000000101110010010101000011110001110110110100010110010011101100001000011010111000010001101000111001110001001110010011000011111010101010001101011000100000101001000101001010100100010101010001100101011100100111011010011000101110010010011110001000010001000011110001001000111011110110000000111101111110011000011111111001011011000110101111101110101000110110011100111001110100011011100000001000011100101010110010000111010111111111111101001100011001100011011000100010111111011111001011101010000101110101010011010110011111011011010110101011110101011110011100111011010011111100111001001011011011110100000011001000101011100010010101111101011111101010100011111100000010111110110110011000010010011001100100101100101110100111011100100000011110000000110011010000100000111001000100111011101011100001111010111001010000101110101011100011111011111101001011100001011000100100111011111110011011110100001011000000011100001101101000000110101111100110001001000111011010110101101101111110011110101110000101001111000011010100000000111000110100111010111011110010101011011010100011011010000101000100110110010010001111100010110111111010000011100101101111101111000101101010100001111111101001110001000110000011000011101101111001111110110000101110100000111110001101001101000011111010101111010000001110111000001100111110100110101000110101110010010001011010001110011001101001101010010100101011110011011100101111011011000011111101111110111010100001100100101001100010010101011100011110101010110011101101110010011011111010101110011100101110001100000111110010101011000101011001111101110111001101100000010010000001100101011110100110001011011000001001001001010100110010110001010000010100010010101101011101100011010101111100001001111111100000000001101101110101010011010000101111100111100010001111010000100011001011101001101110110101110011001001101111101111000100011111000010100011110110111101001001010110001001000010110010100001110101110001111000100010010101101101111110110000011010001101111111011100100001100001001000011000111001101101010101100110101010000110100111010010110111001111111100000000101011011000001000000100111001111000000011111010100110101101000011010011101011000110101000010010101001100101100101101010100101100110001011000010010011111001000100010110000101100011001100001101111110000100010000011011001010011110010010011101001100101001000100111100000000010011100111111011010111011111010111101011100100011101111111011010110110101110011110101100010101001011101111001000011111000101010000001011111100000001010010111101000000110100010110000101001100111101011101000101000000001110101010111001000110001011101010100101011101110111010001000111101001011010000001101100011001110001100101100001011001011101101100011010110100110100001010101010000101100100001111101101000011101000110110000011111011001111111011001010001111001111100010001010101111100111100111001101111111010111000001001110110011010111011010101110101110101000101000100111100110101011110011000101111100001101010101111110101011100011011000110010000111111011111011001011101000100110010000101100101010101100000010100110111011001001110000100001010100001000110011100100011101010011101111011101011111111001110000001111111110111001001110011010110101101010001111011000110001110010001100000011001110011101101010100101010001110101101001101101010110100010101001011101110101101000111111000000110100100111011110011110100010010110000100111111010010000001000101101011110110000110100001010011110111001000001000110110101000001111111001001111111100101101011110101010010111111010011000001100111001000000110010100000000001001011100101101100111101100101110001101000111111100010101110001111000011111000010011101011010010111111000011010000100111001000010011011101100100001010010100111000101101000010101110101010011111101111011101100110011101110110001101010011011010001010010011001110110101001010000101000001001100000111101000011110001000101100100111000110000000011110000000000111010010101111010010001011000011010001000001010011100011000100011000110011000011011001000001100011000101010001001110000111000001110001101110101010001011101101110111001101111100011111101100010001011100101110000100101110111110001011110001001011011000101010001101100010111110000011110111010110000111000111100110100111101001111001100010101011110100110010110000001000111011001111000111000001001001011100111111110101101011010110010110001100110110011110010101000010101001010001001011011001000001110111000101110001011010101000011101101100100001000110011001011011011010011001001100011010001111011011100111100111100001101100101001001111111101111100101011100011000101110100100011101011011011010111001111011000000010011010011111100110100001100001000101110011111101110011001111010110101110111101010010001001101001110101110110011011001100000010000111100001011011101100010000100101110110101101000101110111101111110010110100111110100000100101010010011000000100001000010101101011010111100010001101111101001011010001011100000110011011110100010100001010100011101110000110010101011110011101111100011001110010101000011010101010000111000010101100010001100101101100100001101110001101000110000001100110000111010011000011011010001001101000000100010111100000010001000100011101111100110000001001011100100110011101000110110010000111010111100011111100101011011101101100010101000101001101101011101100111101010000100101000001001111110001000100100101100110001101111110010000010100011011100111111001010111101000000000010010110110010101111010111010100100001011001110100001011100101101101110000011111111101110101110111101100000010101011111110111111110001110110011100000001100011110000100000011011100111111110010010101100101010010111000001011111010111000000110000001010011011100001101100011011001011111011001110111100101010101100010110011101100011100100010100011001111110111011101001101010111000000101000010001001010010111111111111101101100011101111100111110100010010000100001011011111110010010000100101010010111011101010110001110001111001000111101111100101100001010110111100011010111101101110011010000001010101100100001101000100111100100100001110001100111011110000101100101011011011001001010100001100010011001110010111000000010000110110000011110000110110101000001010010100011110100111111000011111011001100011010101001101101011001000101101110000011101011111010001111110010001011100100011110100001010100111110001111110011011000111101100100100101111111011101011111100011110010011011100010000111001010110110100100010001101100100100100100001110000101110110111110101000010110101100011111110010101010010011101111100110010001111000011000000000000000100101110101000001101000111011111001101011000001001100000101001100010100001010101101100111111000101010001000110111011001111111100011101110011100110011100000000110000010100101011110000000100110001101100111001100001001010101101110111011110111001010110100110110111010111100111110111110000110100101110110101011110000111011000101010100100111110110110110110011010111010000100111100100011010111010110111111101000011110001110010111000001101011110101011100100011010010000100011000000001100010011100111010101100101010000010000110011011011011101011001011110101110101100110101011000111101100100010010011011000110110010100101101011000011010000101010010111101110010101011111000000101111110110100100101100100111000110001010100010011111000101001111010011101011110001001111111001101001110111110001110001101000101110110101011100011110110001101001000111111101110011100100110000111100100001010101100111110010101001110100001100001110100001101100111011010110010011010010001011001001001010111110010101100010001111010011111000111011010001110011011010111011011011111001110110000110001111111100011111001001000010011011110110000111010110000011111000101001110000011100000111100100011100010001010110101000100100010101110100001100001011001110001000001111001011010011100000001001101101110000010010111111000011100100100110111110010011010011010101000100101100000001100000001111011000100101010110101010001111000010001100010000110101110100010011000000010000000010111110001110100001000001101111111001000011001011010111000011101100110000101000111001001001001001110000100000010011111000101001011000010110000111011000011001001011110010111110010001111001101001011111000011100100110000001001101111010000010110101011100011011110110100110001010111100110101111110111011000110000110000011100011000110001000111110000000101001101111010011011100011010001001011111101100000110111011111010011111001100100010001100100011001100001010001110010101010010001111011001100011101010111000101010111101101101100011010000111110011001101110001000111001011101010001110100110001011010100010111100010110101110001100110010111111110111100111100110111000010110100111110111001111111011001100011111011111000000010011001110100001011101011100111111101000110011111101110010001110010000011001010001001101110011111000111111000001010101011011111111101101010100101111000100011000000101010010001110111110101101000001100101100000000110110011011000101001001011101000110100110111011101110110000001100011111010110101100001111101010001001011110100001000010000110101010101011011000011110111011110100110010000110000101011010011001110000100011011101010100110110000100010000101100101101010110100110010111010010010010110010000101001111011101110010110001110011010111100101000011001101110101101100001100011101001111101111110010000011111000110100100110000001011111001110001011111000110000001000000101110010101000111000110001100000011111000100110011001101011101010010111010100110101010101101100000111001100100000111101110100001100010110110100111100011001001110110100111100101010011011010010100010110100110010101101010010010110000110001011010011111001010101000100000111001010101000010000100011011011111000000011111100010001110010100111010110110010100010010000010101110100011010101110010001000110100101001101100111101011100010010101100001110110000111111001111100010101010111001110000101011010011111011010101110101100001101100100011000011101001101110001101001000101110110110101110111111111010001010011110000110010001110101011000010001110101100000100111100101001000000010110011100001001111001011010001011101011111101011010011101010011001100011100100110011111111011010011011011110011101100000010011000100011101100001101000011011110111010110010011101001101011011010111000001001011011001100011111001000011001010101010011001010010010000101000000000000001100001011001000111111111001011011011101111011101110000011001100100100100111100010000011101101100011010110011011011011111010011100010101001000001001001101101111110010000011101101110000111010100111101111011101100011001100101101000010101101010110011100110010101110101101001000111110111111000000110010100101011010101010011001000011001011101110111100101000101010000000110111000000001101101100100010011101011100010000011101100000000111111100101111110100011100110101011111000010001011101010111010110001011111000101100101110100110010001000010111011100110100110010010000001111010001110111111111110101110000111101110110010001001111100100010001110001111010000110100010100110100011110110101100111100011101000011100010110101110011001110010101110100000110110001100011000110001111111101001010010100101110101101110110010011110010110110111111101100000001011111110101010011100101001110100110100110011010100101010001100110111110111111100100001110001011111100000111010100011111010100111100100111000000000110100011110000010000010110110000000000011000001000100110011011100000010100100110111001101100000101101100001100000000011110110111011011011101101100100100100011010111010000000000111111100111101011100001000111100110111010001100100100001110000001011011110111011110001010101110111010000101111011110011110110011000101001111100100101101101110110011111010101100100000010011001001101001000111111000100100001111001101111000110000011101000111000111100001110011100001011111110000000011001010111111010011100110011101111001011100111011101011101000001101000111110110000100110101011010010000101010010010111101001011010101001111011101100010101010100111001010000111010011001011000111000100010110011101101010010100000001011001100100001000001011101100111110000101011110011000100100101100101000011010101111100000101110101000101110100011100001111001001010110000110111111110011001000111001011011101110011000001101000100011001001100001000100010101011010110001100110101000110110110111010111101111001100100000111110111111111000011100011001010000001011011110010110100111110110110001101011011000000011010011111110000000011100000111000110011100111111001110110110011111001111001100110010001011101010011101011111100110000111111101110001101011010010110101001000100100011011100011110011101001001101101101011010010111001111101101001101010010010001000001001000110000000100001101010100010111010101110001110000010000001011101111010110001000110001100100011000010101110100011010110010110010001011000010101110000000110110010110001010000000001111000100010101100010011101100110011101000001010110110001010101110101100000000010010001111110000011111000010111000100111000101001100010100100101110001110001111000010011101111010011101001011100000010100101010110111111010000001001001011100110110011010010011000000001100101011010101000101101101000011010011101001110001001110010010100000010001111111110001111100110011111001001011000001010100001000001011111100110011011011101111101110010001100000010100000011101111010010111000100000000101100001100110011110000001110000101101111010101000101100100001010011111100100010010110101100101100000101101101101110110110010111110010100110100100101110010110110001111111010011010100100101100110100001001011010001000011101011101001110100101000111110010010100111001110110001000100100111110100101010101011011001001010110100101101110001011000001000101010111110000110110001111110110100010010011001111110101111010010010111110100101110011101101011001111001111110101001110000110011111101100001100110110100111001000110101111111100110010100001111001001110011011110110111011110100000001011111000100000000000101100111100111001111110000010101111001110010010010100000100000001101111111101000101000001110101010101110111111011101100110100100111110110010011110011000101011010011010111011011010010100000011110010111101111011101011111011101001000000001110000011101000111010000101111111000001100111100011010100001011111101100111110110001111110001011010011110110101110001111111101111111110110000011010001100101010010111001010010101111000001100010101011010000101000010111000001101001101110010001101100011000000101101010111111101110000010010010010100110011000011001111110110111011000101010001110110001011101100010101110010100110101001101001001010010100111100010011101000001100011101100111111001101011100001011110111111010101111101001000000110110111101110010000111010010011011101011101101000011100000000110011010011000100001101101001000001101011000001001000111100001110111011111100111110000011001100100010001111110011001111010011101001100111101000110100100001010010111000001100010000111010110111101101000000001101110101000111001110001000010001011001010110010110111011011001111101111100011101110100100011001110110111100111101101001000010111100000011111110000100110011111001111010011011001110101011111100001111000100100110010100110100000100101000110101111101001010101000100101111011001010101101111101111011011010000100001000011000011010100100111000111011011101110101111100110100010100101111011011010000000110001101100001000111111011011101011000011100100111011111011001000111101111000111011001110111100110111011010101000000010001110100010101110010101001001101100001011011111111110111100110011100100101010101111010111011001111000111000101100101011001111100011100011110110101110011001001100011011100110001011101000100000111110011000000000100111100001101100111010111011111100100111000001010000010110010100111000000101001001111001011100110010011010101000010110000110111100001010111011010101100011010101100011101001011000011111001000111111110100111111110111011010100001110001101000101000010101110000001000101110011100011101101001110011001100011110010001001110100010010000101111010011101011001010010001000111010011001001010110110000011010000011010010000110011110100101000011011111001000000111111000011000101011010000000101000000100111011000011101011001011010111011001101011011010100011011001111110111101101010111000100001011010010011000011010101011100010011110000100011111101110011110011001111110110100011110111010111010001010100111010011110100011000010001000111111000011001011111001110010111010100000111011111101010011001111111101101010100000010110101111011010001011111010101010110011110101010111110111001011111111000111011100111110001000000001010110001001110100110000010101011101000010110110000101111010101011100011010110101100100101000001100100010111110110111100100111010010010110111011110001101110010101001111101101011000101011100001101011110001101000011101011101001001101010101001001100101100101010011101100011010010100111110111111001111010010101001110011111100011001100110101110110101110100010011010010010110101100011111101111001001101110000110110111010101111100100110010001010011001000000000100101010000110110111000001001011010001011101101011001111001111100101111101011100100111000101001000110100010110111111111111110010010001101000101001011110100111001010010111110110011101010011100000001001010010111000010101000101011110101101011111100100010001110111100011100001011001000110100001110000011011111111100001100100101110101101110101110111111000101011110100011100101111001011010011011101100111101011101001001110011000110011011100001111111000011001001001010011001001111101000010010101010000011100111001100011011000110011011101110010110011000110011000101111010100111111011010101111000110010000011111101001101000001100000101010100001110110110000101100110010000010011001101010110111011100001111011101110101111110110100101110011110001111010101010101011100111011010000001100101000110101000111000010101001101101110111001110111110101110110000010001100000101110011101010011100010101100111111101100110101101000010111100001101110100011110001001011111001011100101010101011010111000010100100011011001110010100000110100100011010111001010000101111010011101011110100000011101010011011100011101101000001101011100110010111111110001100010001101011111010111110011011110110101010010010010111000010001011111101011001011010010000111010001010100111010100010110000110000100100001010000110111101101011111101100111010111010010010111111101001110110111100101010100000010100110110110110001111110110110101001111001000101110110110100110010001010011110110111111001100110111011101010111010101101001011101011001000000101111001100111111010000100010111110000010111011100110101011000111100001101000110101101000011000111111001000011110100010100110011011010000100001101101111011110110001010001010001010001010000111101100010010011101110001100100101100110111100001011000110011010011101101001001110110000001010110011110001101100111110011010111110001011100111010111101101011001101111010000011011001110110010101111101000111000001111001001011010110101101011111101111111110000100101111110110011010110010001100010101010010101111101011111011010000100100000111101101110110011110101011010000011000111000010110111100111011111100101001100101101000000100011111011100100010011011100110100100101110101001011001111000000110111001000011101110110000000110101110001011000111010010000010011010010100101101100000101001100000100101011101000011101111101100101001010111110000010111111100111100100110010100101111011010011010000111001101011000010100110100010100110000111000011110101001100000000000010011101110101110111011000101001000010101010001010100101110101001010111010111111010011111011010100010111001001111111101001000110010010110101001010000110011110000100110100101010010001110100100010111010000001001000110011001100010000111100011110100001111000001111000000111110111110000010011000011000101100000101100010100001011011001000001010010011000110000111001101101000111101110001001100101010011011101000011000011010000011111111110110010101001001100001100001010001110101111001001010101101101011100110101100000011111010100011011000011000010001100111110001110010110011000100000100010000110010100011001110011111100110001011010010010100010011110010011001001000111001110110010010111100110110000100011001010000011000111001100011011010100110011111100011000001010110011110100101101110000000110110110111100110100110100110010000011000000000100000100110110111110010101010011010110111100001111000110010110000000100000101101011100111010101001011001001100000111100110011001110000110011100110110100011101001100101101010001011100000001101100011111001100111100011010011111000110001110110011000111100001000101011111001000010111101000101101111010110111111000011010010111001110100101000001101111010001111001110011111101100001010001110101010001110110101101011101011101100110011101110101101001100110010101100000011001111100001011110001100100011001100100000111111001100100110111001111000011000010101000100010100001000001011010011110001010011010101101101101111010101111100001100010001101001111000101000011111011001011101010111111110110000110111001000111111000010110100111011011111110101011000110011110100111101100100010011101100000101101101111101101000101101110100100010011101110010001111010011010000001001000010111111011111110101000100001111011110100100001001000110110110011000100101100001110001101011010110011101000001011100010101101101000101100000101010101000001010001101100100000011001011001111110000101000011010001100111000011100111111000100101001100100011100110111010110110000110010111101011000000100010100001000101101010000110101111101110011000010100101001111100100110111111011000101010110010001110000110010110110010000110001000110101111000010011001100011011101010001111111000011111100110110010100110001001000001111001110110110100011101011100001001101000000111101100100101111011010110000000100011001111001110000010111110011110101101100111010110000110010110111001101001011101010000010111100101011101110110101101010101111011100100001010110111100100010111110010100111111100110111111011011110000011110000010101000010001100001111000011001001110110101110110110011111000100110011010000110100000000001001011100111101110100010010011100111110001000100100001101100000111110010001110010001111101101011011001011100011110100110010000111110010101111110100101100100111000111001110101011100100101010100010111111111011011101000111111011100101101001110000110011011011100110010011001111011111001110010111110110000011010010011001101110110101000011010011101110001101000000110100101010111101011110110110110100000101010110100101011111101000100000011110011000111100111010000100100100000100001000001100110101111000000101111011101111010111011010000011110000010100100101011100001111110001101011111000110011010111111111011110001110011010010111001010100010010011011011001110100011101111010000000011100011101110101111011100100111110101110011001110101001000010011011000000101000111011100100011101010011011101100110100011100100000011000011011010010010000011000011111101001001001101001010110100001011011001110001111000011111101100111000111110101000101000001000110101111010011001000001010000010100001101011010100111011111101000000100111111100010011001010000011000100011000001101111110101100110100000101011010000100100101111101011100000010110000010010100010110000101001011000010000001001101111100001011100011001100010100011100110110011001001011001110100100110110100000110101001110000010111001010111110011111011010000101001010110000000111011101011010001101000000011011001110001000010101101100110010000100010001101110101110011001110110011000111010110000101101100110100111011111010000111101010001010100100101001111000100110000110111000111101011011110111000110001101110101000011110011011111000111001111111101110011000110010110100011001111010010010101100110101000110000111011001000011000110011100111111011000100110001010000010110000111000111010110111111111111010001110111011011111100010101101111010010100001101001111011001011101101110101100001101000000111111110000001000000011001111100100010111100000110011100110011110010001100100111011011001000110110100000110010100100011011111000010011010111011110110110101001010000000001011110010010010000000001000001000000001110101101011111001111011110111011100010111010000001110010101111001010001011011000100010101010011010000111011110110111000110011101101110011101011101010101001100001011111110111110110100111101010001011111000100110011000011110110101010010001100111100110110010000111111011100101001111100001001101000001110011011001010000011010101101011010010001001110111011101001100001010101110110010100000111100010010110110011000101100011101100111111101111000110100001111101100101101100111011001111110010011110111000100110010110010101000010110111111001011101000010110110111110001011011111101100000100010011101101000110111001010000010100001001101000101010001110100101111011101001101101010111000101011110111010111101101000110101100100010100001011000000111101111000101011111111110000000000011101101101010100001000010111111111101100110011010010101110010010101011000101010001011010100010001001010100011011101000001110001011110110101010101110101110110011111110111100111001000100111000011000110111101000001010010011001011110101000100111101000001010001100101110010111101001101100101110001110000010001001111010111011101111111001111110011101110111000001010101101001011010011011111110101000110001111000010010011110011100101111101101001011000010101110110100010010000001100101111010010010011111111100111011110000110010101111011111110101000010111001001111101011000001001111001101010100000010111000011111000000000101111011110111011010101001111100100111101011100111011000010001000000110111100000011001111001001101010001010101011010101110011011011101111001111101110011100001101000011100111111001111100000100011000111101000011111111111001100110010110000100111011101111101101101011001011000110100100111110011001111110010101000111001100101101111011100111110110100010100100111001001100100101010011001010101000000111111010101010101000011110100010101100011111001010111010100111010111110100111001101110001100110010010000100110011110000110010100010101000011001101101010101011111000000011001001010110000001010110110100010101011101000101110101110101001100110110001000111110101001010000001010001001011001001010001011100010000000011100010010010010111100000101111110000100010011101110101000110001111100100001110100010000010101101111100000001111001011101110100000001010101100111111010101001000101101010111111010100000100101100000100110100110010010101100100001000010000011100001111110001101010011011011101110100001101100110101111010100110100111011100000101010011001110011101111100100000110001110111111101010001101110111100001101111001001001010101100101111100011100101100010011101111110010100000101111010011001001000001011001000101010101000010010110000110101011010101001110010101010111100001011001101010100101101100000110101011000001000111010111101000101010111011000010001000110001110010010111000100000110001001100000000111011001001001101111100101000001001000101110000110100100010101010001000011101101010011111111110100010000001101011011000011001111100011111110001011011011110110110010011100110111110000000000001110011010111101111000011011110100101101111100011010000101001010010010110101011011011100100100110101011110001111011101000010111011001011101111011100011001001111111110100110100000110110110010100110000010001010111010110001011010100011001000010001001000000100111000100110110000011100011111000110010000100101101100111101101010001111111110000011111001111101011001111000011100001000100110000100011001001011000001010010011101001010101011111010010110000101011000111101110101100011111101110110100001011000110111001101110010111110011111101111101010011000100101110010000111111001011010100001100010111010010101101001100001111001010010100101010000011010100110110010111110001010100110001011011000010011111111111101011100000110111010011010000111111101101100100010111011111110101101100001000001010101101000010101010010001101110101111010110010111100001110110001110011101010011110010100100010100110010011010100100111011001111011011100000011011110001011010001110111001100101101110111111011110010101000001011010010001110010011001100110010011010111011000101100010101001101111100101011101011001110001110011001101111001110011100001101010001100111101101000110010011010111000111000010001101111101001111011011010011001100010010011000000101001001011110000001100000010001100000110011010110011100111110111110111110011101000001111111001101001010101010101000011000011010000110011101110111010100100100110010011111010001111010110001100100000100011000111011110100110110011010101011001111010111010101100010110100100110000010000110011000011110111100011010111100011010000000101101101010110101000001111011111101010111011100101011010110011111110010000111011010010010111110100011100101010010011011101010001111110011101010011110001110011111111001011001001010001111100101000000111100010011010110111000010100001011010000100000100111111100110101011001010110011011111110100011001000000101011110111001101100010100010000110101001101000000100010110011111010011111000101011100000111001000110111001111111000101000101100100010010100101111000001000100100011111000111010001010110010011111001110110000001011001110000111001001001011011001100100011101100110001010000011110100000010010001100011101001100100100111010001011111100110011100011010000000010010010011101110100000000001000000011010010100111101110001000000111100001110111111110010010101101101010110100110111001011100001000100010110111000111010100010110100011000010010010011100100000110100010000010100011101010101010111110101001000101111000101010110110111010011101100000100001011000000111100011101101010101101010100101000010000001000010000001001010101111100101111010101101110100001111110101010011010101011011000111010011000000000100000001111001110101101010111010000000000000011100010110101100001011001010010111010011011110011101010101101001111001011101010101000011001010001011101111011001100110101100110001000000111110100010111110000111010011101100010101100011000110100000010010110110000011010001101110001100011110101010100010111001100010100011001001010100100100000001100000110100011111011011010100101000111010000001111110000010001011110011101011000011111010111110000001111011001100111110001011100011011100110110010101101111001100011001000010110101110000111011110100000100101100010010001101001001111111111010001110000000010101010101101011000110010111110110010010111110001111001011100111111101100000100000111110010001000101111110101101111110010010110110001111101011110110000111111010110101001110011110010001000000101000010001110011100011001111101000000001001011111010010110100111101100111101011011100010011101001001101101011011111111001001110111111011011101011010100001101111111101100000101001011000001100110110001011111111111110100010101011111010010111001101001010011010001101011000110100110101010011110001111111100011110010011001001100110001000011100110010011111101111000110111011100110010011101110101100100010110011011011001100010110010000100010001011000010111110110001111011111001011010111111000011111000010101110101000010000001000011110110100100001001000000101010100010001000011101000000101101001011001000110000011101100000000101000101100101100111100010010011100101010101001010000100101101101110001011101100111011100100101101000011000111001110001010011110011111101011100111110010011001110001010011100101010001011111000100100111100011010111100100110011010001100000010110001011010111111010111110110100101111111001001100100000101100001001000110011100111011010001100011100111111001111111010101010001011100000001110011110111010101100110000110100011011101010101011010011010001000110111001000010100100110100010100111110100111000000001111010000111001000000110110000000111001010010110101001001001010110010010110010111110011000111011011111000110001111000010000010010011010110010110000011110100111101101001010000000000100010010100101010000101010101111001011001100110010001101110010110110110001110001100110100010011010100110111010100011111110011110111100000010100101111010101010010110000111101110111001011110001111011110001110000011111111010101000101110010101111100001101111111110001110101100100100001010001010110101100110111100101100110000110011000111011111010110100000101000010011100000011000011011101000110001110100101000101101111111011101110100000101010010001111000110101001001010101001110010001011100011111101011111110011100001000111110000101001100000000110101011100001010000110010000110011000001010010001101100011011110111101111000010110100011011001110010010011001011110111111000010011111011011111010001011010101111110101101001110111100000101011000111111010011000000000000001000110111001000010011001100110101111110111010101101111100011000001110001101110011101110001000111011010000101110010110100001110010101000001001111100010001100001100001011110001001101110101001111000111101000101111110101011000101100010110100011011011001000011111010101010101111011000001111011111111001111101000010101000111101110010011111011010100111010010010100001101010110000010000011111111110011010101011101011001011010101101010010111010110011010000110011110100101001011111111001100010000000001000110011111110100011100110010011100110100010010111101110000111101010000111000110001101011101111000001111101001000010011011110010001100110000001100001100000001001000001010000000011000100011101001100011100110011010000000100011111000000101111110000110111110011001001101001010010010010110010000111011010001101000110010001000101100111011110011011010111111110011100001101100100100101011111111111000000000000011111000100000100010000110111001101100010101110100111011011101101110011101111101001011100100110010000110100101010111001110001011010101001010111110111001111101011011111101111000100000000100110110110110101100100000101110000000110000110000001011101010000101100101000001000011000110100000000010001101111110110001110100101001010100111010010000101010110001110011001000110111010001011001110010111001111100101010110100010110101011000010001000010111000100100001011110101011001011101000110001011001000100111000100110101101011101111100111011110010100001111011000010010101110101001011001110001111001110111001000101101001111110000100110010100110100100000010001100100001111000001000000110101100101001110000000110010011011000100100001000110101011100001101111001110001001001100101110100100001011100110101100100010010111111010110101000001100110110000000010001111001000011110001110010010110101110111010100010001100100100010110011110010000001100010001010010000100000011000111001110010110101000100111000011001001110101100000111101010010100011110010010100010111100111011010101001010010110011010110111010011111010010100011101110011000101111000011101111110101001011000101000000111011101000110011011011001100000110110110111101010000000000011011011010100110111101010110111011110001110111001001000011110000001101010101101110001110111101001010010101001010111010100000010110101000001011111000001011110100101101101000000101111101100011010110000001111001011111010111110101101101001000001001101101101011100111001011000001101110000001001111110111000010000111100000010011001011001100001000011101011000001001000111001000010001000010101001010000000100111110110001000111101000011100000000011001000000011010100000111101001000011000000000101100100001110111011001001110101010010100110111000010110111100010111000101111001101000000100110111110110110010100010010101011000011010111101111111110101101111100011001010101101000010100011101101110100101100011111100101110100010010000100000101100010110111110000111010011111001101111111111111011101011101011011001101011101110111000001011000101100101001001101001011011000010001011100011110011010101100100111010000111100010101000001011111001101100111110100001000111101100100001111100101111000111110110011111101001011000011001100110110101110011000101111010100111000010101111000111000010110101101111001001110011100000010011110111101101110000111101111010001011111111100001010101010110111101101101001111001000101101011101001001001001011101000001001010111011010010110101110000011001000011111000011011010011100111010000010011100000100101111111000100011010110011100000110000100110100100000011100010000010010001111010000100110000001000101010111010100111111100101000010000100100011100011101101101111111111001110001101000001100111010111100111110111010110011111011011010111111010000100001010111000100111010110111001011110100110001000101000101111010111011101100111100010010100001010001011110010001010000010110110111011111010100011000001110101011000111110010000110110001100101001101111010101101100111010101011101000001111001100000010111110011100000000001100101111011100111011001111101110101011000110010000011110011011000101011100000011001011010110110111100001000010011110110110001011000111110011010101001111001000000110101101110000011101001001001111111000101101110000011010110110110110000111100100101000000101000001101110100001111011010011101100001110111011001000110110101100100010110000111101101101110010010101100010101001110111100001100111000100010001000001110100010000110010011110111110110101110001101010010001110100110010101101011010001110000110000000010111001011110111111100100011000001110111111010011011000001011011111101000001111110010011100011100110110101110110011111101101001101000100011111111110100100111001010100101100110101010111011010100110111111011101111010111111010110001010100001011011110101110001111101011111000010001001110000001110100110101011000101101000011000100111111101011100110001001010111010010001110110001101010101001010011111001010011000101010010000011110010111100101101100100100010001000010000000100001111100011110100111000001000001110110111111101110010110101001111000101110011100111000011100011010011011010010000110100101010000111000011111011010000101111111010100000101101011010100000110101000010000100110101111100100011101101010011110000101011011010101100100111100000100011111001000110111011000100110101111101111100100001101101111100001110000100001100010011101000110011011001000111111111000101000010001101111110001101110111000110001111010001100110000010100001001110010100111010100011111000101111101011100000011100001001000000100100101000011000101111111100000101010011101001000010101000111001000101000000000011001010000101111110110010111010101111101100100100011010000111101010100100100011101011010001111011111101011011110011011100100010110001001000111110010111110000001010111111111011110000101110110101101010011110001001101110111000110011111010001110100111110111000011010110100010110110010111101010111000001111111111010100101011001001011110110000000111011110001111110001000110000111010011010010101100110110100010001010010110100010100000101110101000000100010101010111011100111011100011001011111011001111011011011101000110110011101111100000001001101001011100010001111111101011000011010101110101100010111100110010010011011111101011011111010100010011100011001110011000110010001101101100110011011100000110010001111000010110111001011010111001010111001101111110011001011101110000100101001011100110111100110000001000100111100011001000010110111110111100101001111001010101001010001001110111010001111001011000110010001101011001011011000110110110110111001100111011110011000001001000011010011100110110010001101100001100000010000101101000100110001001000001001001010000110001000001111111011111101010010100001000001101001110111010011110110101010100110111100000010000101000011110000101000010111001110110111110100010110101010010001000100111011000000011101111111010010001111101101111011110111110111000110110000110100010101001110101101110000001010000001101100111101110000010010101111110110010011100100010101010101011101000000011000111010000101011001000011010010011110010111101000011001011001000110100111110110101011010000110000111111011001110001001111101101001011011011011010001110100110001111100011110001011001000111110100010010010100011011101111110100010110011101101101110001101111111111100000100101001100101000100101001101000000100001111100000111110011111110010000101111011100001101101101010010001111010001101110000001100111011110101100010001000011111001001001010101001001100110111010011101001110100100101011111001001111110101110101111001011000001100000010000000100011011010010000101101011101011011000011110100111110111011100111100001010000010100100000101111110011110111000001010001011111101110111000000010101000001010010111000100101010011010100001001010001011111111101111011011010110000010001010001111010110001000100111011110101010110011001000000100111100011001101100110100100110011101110011001000010001011001001111101100010000111010110001101001011100101010001001101101100101011111110011011110111011010100110010011100100101000010011110100011111110000011111101101011110000001110101110010110011100100000110010001000001101101101010001010010110010010100111110100110011101011101100000010110001111101101010101110100010110101000011011100011100010001001111111111001111101011111001101101100100010101010001111110110100100110000111101001001111111110111011111110110010101000100111011000010001111001000000000110101000110000111110111110000110001101010110111000100110100100000000000110100101010110101110111110011011110010100000011010001111110011111111001001011001010010100110011001001111110011010010000111011111100001011011110100100111011010010001000010110100101101111100000001011101110001110000000101100010000001111000100100100011110000010111010101000000101110000000001001011011111011011111011010010001010000010011001111011001111100001111110101001010111000000001011010101001010000000011100010110111010110000100110111010001100010000001001011111010110011100001010000101110001000011101110000000110001010100110000000100011101000010011010110011111111010111000001010100100101111000011010001100111001011010101101011110100110110010100110001011101010100001011100110110101010001100110010000100011010011110100001011000111000101111111111101011001110011001000100111111001010100101001000100110100111010010010001011101000010010011101100111101101100010101011011111001110101000001010001010110101011001111011101110111000101100100001110101100110111011110000111100100111000011111010110010101000010101011000001000111010011000110010001110111100111100000110001110000101010010011001110111001010010011010111100010110100000010111110001011001100111000110001101011111110011111010111011111001000010001010110011000001011111000010101010100001110011111011100110111010001010111101010100101101110011110001101100101110111111110111101010001010000101101011000111010000110011101011000011000011001100011000001001011110111001100001001110101001111111111111010111011110001011100101101010111101011101010010001000111000011011101001000111000011011001001111110101011100100011010110111111000111111000001100100001010111010101011000111001110111100001110010001111010000011110100101011001000111101110110101100000100010111011011001001111000110010001010010101111110000000011001001110001111111110100110111101101101010011111010111011101111010100000001100001100111100011010110111101100101011000001111101000111000111011111111010001010101000001111001011000010011011001011010001101111001101010110010000011100100111111000101001100001011101110000101000110011111000000001011011010110010111101111110000110010011000011010001110101111011100110110001100000110001011011100000011100100001111110101100100111011101100001010110110010011000100110100101101000001001100000100111000110110101100011000100101110010001010001100011010010010001110011110010000101111101010000111010110011000001010111001001101110100000010111011101101010110011010100000001011111101100000010010111011010000000101010110001001110111010001110011010000100011101011110111001000001110101011101000010000010010110000110111100000100110101101001110011011001101110011010111001100100101111000100001000110011011111111011001111011001100100000100000100110000111001001101100110011010000111011111000010110110101001011111101000001111111110010111101010111111111010110000010111110111010000110011110101110100001110011101010111001000011101111111101101011101010100111001110010010100010010010010011000010010001110011010101100110101010011110011111010111011110011111010011110100011011001001111100011000000001011110000100111101000000001000011011100111000011011000100010101011011100000100011111110110010101001101100100110011001010010011010011100011011110101001011001001111001101010011100111111111010000111110101001110010001110011111100101110110111110001011100010110110010011001010110001101111000101100110011101101110111000110101011111101110101100011100100000100100011000100110111100010110011111011101001100110000001111011011101001000001001101100110011011001001100011111001000100011110011101000110000000100101110011011011101010101111100101011010110000100111001010000100000111111011010101111010011011011101011100001000111101000111011000111000110011010001000001001100001101011001010001001011010000111010001101111000000110000011101100100101111100100101101101001011101010100010110000010100001100011011101000100110110100110110010101011111010100110101010011000011101110011011110010001111000110001100001100011101000000101111011001101100100100100100011111010011100010100101100001001101110001110111001001111011011000111000111111000110001101000011000100101000110100010000010101110011110000011010110110010111011011010000111111000101001010111010001010000111001001001010111000110000111011010000111010010111011010000001111011011001010111001110110110110101000010000100100101010000010101111010001100100100110101001101101111111011000001001101101010110000010100010010111110111101001111111000000011001011110111001011100001011110100100010001110011111011001111000111011101110110010001100011101001111010111100100000100011010101000000100111101110101111001001110111001111111100001100110010101110000110010100001111110001101110111011010000101110100001011001011010001101010001000101001011011111000110101000000101111110100100001110110100101111010010011001000011110111110010010110101101101001010001111011011100011101001000010110000010010010000011010101101100000000010100000110001111111101100011011100010001001010100011011100101101000100100100101111110111110011001111110011111001110001110011101101011100001000111011101110011000111000001011001011000110011000101111101001111001111111110111000001111110011001111100100111011001100100000011010100011010100101011001001101111010011001100110001110001110101111100000001010010101010001001100010101011001111011110100111010000111100010001000011011101010010101100010010010111101111010111000100010110101111011000110100000010110101100011000010111100011001101110110111010010101111101111011011100111101001010010110110101000010110110000100111110110001000110001110110101110110110101111011010011111011100110000010010100111011101100011110101001000110111010100101100000110111000110010101110010111000101111111100011000101000000100001101111111010101110110010111001100100011011100000111011110010110100010001101110100101001011000110110101110101000001000100101111101010010101101001010101001001011100010110111001111011000100010101001001011011100001010010110101001010001011101101100010110010011000111000110101000011010010101100000100010100100010011010110001111001011010100100111001001101110001000011011001101010101110000101000101011110010000011110110111001010110111110100011111100111000110001000001111111101010001101010101011001001100010001111010011101000011101111101111110111011010001011001011010011111110101100010110011000010010011100001111011011001011111001010001001011000001100001101111010000010111001101001110010010010100110011010101101111001010100111111011001111110110011011100101000111100110000000011100110110001100001011010010100001011100111000100101000100100000100111111111001100100011010101001101011110001100100110110101110011000001111000101010101000101101000101110010001111000100110010110111111101111001110001110001001000011100000110011011111100101011101010111000110111010110001011111100110110110110100111110110010010000011101000110111010001101011010000111000100101110101111000000001101100111101101001011001011011010101101101111000101000010001010011001011111001000000001010100011111011100111100011011100001010010001100010001100010011101110011110000110110111111100101011101000010011000101100001011001001100011011110000101100101100101110010010011010100111101111010010010001111010111110110010100111101111111111100001010000001111110011000011001001010111001101100101000010101101110111011101001101100111000011011011001011110010000111100100100001110110001110001100101011100001010110011000000110011101100010101000111111000010110010110110110001000100111011011000110110000111111000011110001001100101010101010101111100000001100010011010001001101110011110100011110010101110001001101101010110110101011000110110101101100110100001001010111110000110000110011101011000001101100001000011100101000001111111010010100110010000111011110001011010110100111011011011001111010111110100010110001001010100101110011110001111111100000111101110100101101100010100010101001110010000010010111010011001100010001010001010110100001110111111111110101101110001010011110000010101110100110101010010000111010100101101000111101101100100000010001101110010001000110111111100011011001000100011110001010011001110101111011110000100100111001111101111110111110000101000110001011000001000110100001011101101100101111111001111011010111111110001111010010100010100101110110110011011110010000000000010100011001111011111010011111000000100110111101100011110010001110011110010101000110001110001001000110001110111101011110010001100010011011110101001001100001001011100000101000010100111101000101101000110101001100001001111010101011111000111111111100101001010111000011001000001111001001011000111011011011101101010011111101010010010000010111000110001101010111110101010101110111110100010011110011110100111000100010111000111111001111101011010101001101000011110001000011110010011110110010000100000111111100011101111111001111000000101010100001111000101011100000100110001011110101011110001110010000010011001100001000011001010001001111010101101110011010111011111110010000000111110011010010101111100010010010010110110010001001011011011110011111000111000000010001001010010111101011001100100010010000000001011000010111100111011011101110110010110100100110100101110111010101011111101001001010000001010100111101001001001001110011101001000110010000110100000100011010010011100010000010101011010101100110001011011011010011100101010110110011111110110011001110111111010010101101101010010001110011111011000111101101011101100101110101001001001010000000011111100011100111101101001010000011100110001110101111011001100101110110101000000010010011111111000000011010010110011110001100101001011110110100100101110101001101000101001011001100101111000110101111101000110010010011101110101000001111010011010000010100001010110111111000000101111111001011010101111101101000100011111111110111100000100101011111010001011010110101100110011110111100010101101000101010010000011010110001111111101111011110101110101001011100100011100000010011001111010000000110000001100010000010101000001100000010110011001000011011101010100100100110010100011001111110000100101011001111001000110011010001110010100011110011011111111100011010111010111100110010010111110101111001111000010000100011010110111001110000111011100110111111011100110111000010000100010000101100111001111100010001100111100100010011101000010110110001100100010100000000011000101011010111110110001110000111111000001001010011100101010110000001111110101010010000110101110111101110011011010001101011111001101011010001010111000101001011111110111001001001000110011101010101101010011111001101000110111100111101001000010010010110001001001010000011100101111101010010111101100001011000101000001101001001111110100100101001110110001000111100110111111011000101111111110001011110100000110000100101101100010100110011110111110100101000010100100011011011010001000011110000011111111000001001110100000111001110101100000110101000011111100111101111100100011110010110001001000111010100100110000010000001000111101001010000111101101010010100001000000001010100010100001011010010100001111010001101011100100111000101111100110000111110100011100101110011101110101111011000100111011111010001001011101111101011111010001000001100000011010110000010101010101111011010101111110110100100111010101011000111101101110000001111101011110100111010010010000100010011010011011101111101001111100000100110110100000011011000011001010100000001110100101110100000110100010110110101111110000110111000011110011001111110100101100101000001000100101110111010000100110100001010001010000110011010011100111010111000011000001110101001001010011101110000000110100101101101110011011111001000110010000101001011111000110001110110011110110011000000101010001100110000000010100001110000011000100100000011001011101000100010101001010010000011110101100111000010110001111100111000010011010101111001110101001111111000001001101111101000101011010110001100001011001110001101100110101010110010011111100011101100001110000010011111100100110001011000101110000101100000101100110001100001000111000111100111110100000001110101010011011010011110100111110101110010101100110111000011100001000001100101011000110010101101001011010001011100011101000100110001111101011101000110110110111010011101111100010001110111100011010111000000101011110100111100101010011000001011001011001100011001111011010011100011001001010001110010001101100101000000001011101101101001010101111010100110011111000011010000110010100000000001111110000000011010010011011000110010110000010100110100011000100001010111000101001011000001000110100101011001011000101011011000001111011000111011001010010100100011011000100110011000110010111101001110110011001100100101101111010010011111011110101100010011111110110111010010001100011001100000011111111011110111001001110110010100110011111100110011101010100011001011010100111111110100010000001111000100110001011101011001111011000101100011000010001010001000111100010000101111110001101000111010001111100100011000101000101100001001110100010001110110101010110010010000100110010110100001010110010010111000010110000011111011101110101000101011110001010100111110101100010010101111101110111100001101101001100000100110011100101001110011100100111100110011011000110001001100101101100001101010011100011101000111001000000100000011110110011001000011110110100111100110001011001011011010110011110000111000100000111101000110100111111001101110100110111100111100101010010111001111010110101000001000110010011011011001111111110010011100110110101010100000000011100010001110111111000111011111110100001110001100110111110001010111010010011011001100011110010101100001100010111101001101101110100001111100011101000000101100111001000010100100110110111011011010101001010011010000111000000111111010101100101000010111100011001110010100001100101011101000101011011010000010100101110000000110010010101111110010100110100010001101001010001010101100011110000110111110111101010110101001001010111100110000111111000100110000100001010010010001101100010110001110101000001111100010010010110011001111011011001101110101101111011110010110101001100111000001011000111010101000110110101110111100101100100111001001110001111110100010110111101001101110110001111010111110010101111001000111001011011010001110110100000110000011100111110000100100001001101110100100110001011011100101010010100011011010011101110010001111000111100100000010111111011010101000100111110011001111001001101100101110100100100111001001001100011110001000010001011011100111011110111001110010000100000001000100100011010011001110011011110111111001110011000010100010011001011010011101011111000111010010111100000000110001100000111000010011111111000101000110011110011010010000000101001001001000010110100110100111100111111000111000111011101100111011110101010010011011111111100111101010110100000101010000100110011000100001100110000110101101100101001011001000100100010110110100000101000110111000000001000001001111001011010010010110111000100110010000010101100010111111101101110100000101100101001111011110001101011001110000000101000101110110011000101100011101000000110100010101000000101001010011101100111011010111101010011001100110001110000111001100011000111001101000010110000111001110100100000001110000001001100010011111101100000111101100000000001100101101110001000011101101111010100110011100010000110011101011010100000101110001010001100111011011101011011111110111101110010101001010100010111110001111111000001101001010100000100111101100010110011110110101111011011111100001011101001001110001000101000110011110100011100011111001001100001001011000011001111111001011100110011110101111010101111111001000110001001000011110100110110001110000100010001111101111000000011101000101101010111000101101111001000010111000100100111100011100101100001000010100110101000000100001010010111111100011001000001010000011100110100101011011101001100001010100011011100101000010100100000001000101000101000100000101110011000110010110010000001101011100110110000011010011010110001111110111111110011101111000010101000111001110111100110111111001000100110011111111011011011001010111100001001011000011001010011010110111111110111001110111001010011110100100110101100010111111011111001101100000010011110101000001000111010110100111111010010100111111111000001101010110000101010111001011101100010110011111011001101111101100000100011100000111111101010011011001000000100100000001000101011101011101111110100111111100001111000100100001101111111111001010011001110101001100010001100100111010100011101100011001100110001101111000010000111011111011000011011010111110111000000010001111001100101110000101011011001101000010110011010001000011000000101111011111010110000111001001000000111000111100011110010010100110011100000011110100010001001001100010001001111110010010010000101100011011001011010111100000110001101101001100111110111100001000010011010000010000101110111100010000111010010111111111110100011010101010111001001010111000001101010001010101010101010011010011111000000111011101100001000110100111111011001010001110001000111100100011000000100111111001011110010111111001100110001000101001000001110110011100100101110111001010110010100011111011000011010101001000101101000111001111101001000000010010000000011001001111011001010001110000010000010111110111100101111111011101010010000110010100011110001100110111000100010010111001110001010000100110110100010100000100010101101011100111100010011000001101001010001101100101010000011100110000011011001110101010111110011110011011010000000101010010001101010100001110001101110000110011100000011000111000010011111010100110110001111010101011110101111100101100100100100111010111101001111101101100110011000010111101011000010010110111111111010111111010010100101011000011100110110001011011100101010001110001000010010111010100111110000100001010000001000110110000101100000001110010010001101001100000001000110001010010111100011000100011110001111011110100011100010101001101001000001011110010110001000110011011101111101111111010100101111001111001011111001000001010001111101101111001111011010001000000110001110010110110110111011011110000101100001011110110100000111101001000110101000100101011101001111100001000011110110110000011111111110101010101110000011011001000011001110100101100001001011000001010011111101110000100101001010100100111001110111111110110001000100110110011000011011000011110010011101010101010011000100111001010100001111010111111000111001011010000111100000110010001110110011010100010000110110000011000111001000100010011011100010010101110111011110111110100110010100101101010000001110101111101111111111011001011011111110011101110111010101010111000010110111000100001010111010101001111000001110010111001010101110000001010100110011001101011101100010000000001100110010101010111101100100010110110111000110010001010111110001110001010100100011011100101011110100000011010011110001010101010001010111101101100100000100111010101010001011010011011101000100010001001000001001011111101000010010010011001101010101101101011010001010101010011000111101000011101010011010101000010101010010010000010111100011001011111110011000110111010110000111111110110101111000010011000010110001100011101110000101101101100001011001010001001011001001010001000001001001100101000101100111111011110111111000111111110001011011110111010111100110100111000111101111100010001100000110010101101110101001111111011000010100000001000001110110011110010110101110000001010011100001000011001011001000010111001000110110110000000010011000001000010010001110011111000010101100110101000011000100100010010000001101100111011011010001110110000111000001011001111100001001110001100111010000110001111101110011000010011000001010011110001001101111000010111111001001100001111101101111100110000110011001110001010001001110101011010100010111111101111111010100010111000010010101111100010010001110101101001011101010111011101001001100011101000110000101010111000101000101100011111010110111001111100000111111101111011000100011010010001000011101101011100111100101000101111101101100010101111000001001100101000000101100010101011001011100110101011100101111101000111110001101011111110000110110001101110100000110111110001001010010001001101011110001001101001000001010010011001011000011110000101011001100101011110011011010001100011110100010100010101011010010101100011001110000001101011010001111001100100010101101000111001001100010100000110011101000100101101101100010001110000100010011010101010111001101000000111100101000011111000001001100100100111000010110100000010011001010101100111001010001010111110001010110101111010000100001001100111100000010111000110011110111101100100010101000000001010010101110001110010001000110001111000001100111001100011111001011110111001101000000000001111100111000001010010010111000101100110111011100111000010011001000001111000010110000110000100000111101100000000101100001110010110100010001100011100110100111011111111100010100110011100011001100011011010001111110011110110100010001000010011101100011111100110000100000010001010000000011100101010110110010001110010011110111110100110010111111111001100101101101000100001100100110110010000010001101100000010100111111111100011010011010111100111011001100111101010110001001110011111110100110011000000111011111101011111110000111100100011110000101000101111110111011101111010111011011100110101100111011001001001011000111001100111110010100000111000111111111000011100000010000000101001111111001001011001101011011011110010011010001011101011010110101100011000100100000011101000111010010011011011100000111110010010010000000011110111110001000001101010111111000011011011001111110111010111111000110110100100111010000111111010000001111100010001101110000111100000111011010110110011000011000000011100011011011001110001111111111101111111001011000101011011011110000001010010110110010000010000111100001011001000111011000101110011010010101000111000000010011101100101101011100110111010001001011101111100100001111000110100100001011110111111110111001100101001010111011100100100101010101110110100100110001000011011100100101111010101111001110111100110000100110110001110001110111111101011111110100111111101001010000110001111100100110011011110000001100011110011110100011100001101100101011111101111001110001000001011010111100111010101100001100010111101010001110000011100110001001000010111101010000010000010111011011110011101100001000110110001010101110011110001000100100100100101100001000001010011011011010111011011010100111000001011011110111110111010100111000110001111110110111110000101000000101110011100100100110010001110100111001010011101111101101101110001100001100011010100100000011100000111011011111001111110011000110111100000010100011010001011101101110010011010011011101110110100011111111000010000000111001000101000000000100101010100000111011110111010011010111101111110101010011111011111111110101100011101000000111100011110000100100010000010000100101111001000010011001101110110010011011001001001011011110110001010010100000111011100111010011100011010011100110110010111101001001010011110101011110101101001111010110000100101010010001100111100101000101010000110000011010101100111000001010000001010101011000000101100110100010010010111001100110111000001010100110001010010001100110111011101010011000001000100001100111011110000011101011011011111000101111101101010010111100111001111010110000100111110111000100101111100100011101111000001101010100000100011010000111001000100010100001011011100100111011010010000110100111101011111110010101101110010000100101100101001101100111101001001110001101101001001010100101100010000000101010010111001100111000101001001101101110001101111101001111101100101111111101101011111111000001100000011011001010110110101100101101111110000110110010100110011000001110110111100011001001111110010000101000101001010100010001101011101000001111100110100110111001111001001100110101011100111100011111101100000101111001001000101111111111011101110111010100110011011011101100100010001101111100101010001001110010000011011100011100110101101111010110110001010111101101010101111110010100111110001100011100000110110100111111011110111111010001111010101011110100111000101100001110010101011010101001110000011110010101011011010001101110010100100000010101000010011011010110000001100100001000110001110001010000000110011100011111011001010011011000101100001110101110000011101101111101110010101110001011011111001000010001011001110110100100011011010111110110110100100110011101000011010101101110110100011110110100001010100101111101110111011110000001111000111101101000100010100110011101111100100001101000010111000001100010011110101111110100100111111111000010011001000110111111001101011000101110110011110000010110111010000101110010001001001001110010001011100000001110011010010111111001101001000100111100001011110101111110000111100001001011000110010010111100000000010001100010110110100011110001111011101101110011011100100111100110001110110101011111101011000001011101010001110111110100100110100001111110100000110001111001110111111010111101100111100111110110010111001111010000011011110111010100101011001110011001101001011101110000011101000010110010110100100110111101000001101111011010100110000011010110001001001001010101001001100001000100100000100010000001001010011110001111101000010110010010011111110111011110100111011101001111010111011100011011101011110101110000101001100101001111101001111001000101010011001000111011001100001111011000000011010101011000000001010110111111010110000111111000011001100001010000011111011100110100101101010000000010010111001011011001000110001101001011000001011011010010100000101111010000110011001100001010111111011101100111101100011100111001001101110000110100100101011100011110011001110110110111011001001000111100100101011101101111010111000100101110010011001010111000100000100000010110001101110111010100010111110001001011010110011100010110010100111000010011110001100111011110011011010010111010100111101000111010111100110001011100100111101111011001010010001110011010101001110000100110010000011101000010000110110111110110010011000110000111110111100010010001010001010100001011000001110001110110101001100100101001101001101111100001000110000010011001001001101101111110101100100100010101110000111100011110001100100011010100011101111111100101010100011001000100111101101010000010011110110000110111001011110110101111010100110101111011010011001100001101111000000000001111001110011100011110000100011001010100001001011000110001011010011011111000000001010000111101001110101110111011100001100010101011001100101111010011110111000000010111010001110100111101110011000110111001101100010100101100100000100010010110000010011111111111101001010101111010000100011100101000011111010000100000111011001010110100001001000100011101111111001101111010101010111111110101011101011011010100110001111111000111110110110101100100110011000011110010111110110100111111011111010011110100100001001011110001001101100101001000101000010000011100110011101011111001101110001101110101010000101110100110100111010111010000111000111110111110101110111111010101001011100101110111000010010110011010111101111010000011011110000110000110010001000000101011011101111000110010000110100101010000100000010111010111110110100000101100000111000110110000110111111100101111000001110011101000111100101110001101001111000010010110101001001000001011011000110011110111111001110100010100001100110101110100001011101010101101010101000101001100000111000011011000001101101001110001010001100011100100001000011101101000001100011001001010100001111011110110111010110010000101101000111101101000000100011001110001010111011110101010111100011010000100011101011000100000000011000010001010100001101111000101000010111001011000010011010001111101100110100000001011110101110100010100100010110011010011100101111010111110100000010100010010111010111111111110111011011110001010010001000111001010110010111101100110010101101001111010111000011111011011110010001001011111010010111011010101000010100010101110110101110110110000101010111010011111011100100101100011101111001010011001011000010101001000111010101111001111000011110000011000000101000101001011011110100010111110000010010010010100010111010010000110011110011100100100101110000010101010101011101110000110111011010011000110000011001101110000110010000111011100001000010100110100001101110010001001110101011000101010001000001100101110011011110011101001111110111100101011110001110010111011010100101110001111101011011011110010001100000110100000101010010001111101101101001000111000011010000110101101110100011101101101010110010111101010011000110111011111010111010011010110001110111000011001010001010001100000100101010100100011000001110011100011000011100100011100011011100111110010100010011110101010001010101100011011101100000100101101110001110001001111001100111001000000100101110110110000111000100100110111100011001110110000100001110110111111001110111010000111000101101111110001101001001111011110110101011001011010110101000001100101011000010011100110101001011111101011000101100100010011111000010011110000010001100001100001110100110101000101010011110011111100110000101010000110001100101000000001100100100111010101100010010100100100101001000000110100111001000111011010101100001010100111010110011010110110110100011100111110011010100100111000010011111111100101001010101101111000100011000011101100101001001000100011001101110101000011000111101001010001100111101111010111001000000000001001110110011100010100000111010100101001011010100101011110110001110110111001000010111100100000111000000101110110111111110010011101001011110110111111011000111111111000101101101100101110011110011110000011111001101101011010101000111110011001100110001001111101001111110100110101100001000110011111010010111101100101100001110000010111000111000111100000111011110000101111110001110001001011000010000101010000001010100001110001010010011000000010100110010011011010010101011000110001101111011010110111001000001110110001001010011111110110110000011011011101110100011110011111001111110110110011110111111011100010011101100110100000110100001010101110111011011110110010010111100001001010011010111100111011110101011110110001101111010000011111010011100101001010100010101100010111001111011011100110100110101110100110000001111110101101011100001001100101110100101001101111010001101011111111100000010001101011100000111001101000001100110100010100101100000100011100110101011110000001100100010011011000100011010110000010110011010000010110101010001111000000110011001111000010100101111011011011110101111111101010100100100001000001001000010010111010000000001010110100011100011011000011011110101110011111010100010001011000110001110011110110111010001011100011101010010010101000101100101111101011011111100011011001001101110000000110111101100111111011000100010011011101001101010100110110101100111000011001010101100101011011001000010000000001000000000001101011010100001000001001100001100100110111100101111011001000101001000000110010110011011100111110010111000110110010100010111001011101100101010110001100101001001110001100111010101011000111010100001100000101000110001111110100110011100011100010100000000111001110010001000111100001101011000111000010011000010111000101010111110011110111111001010010000110000100001001100000011000110100000011010100101111100010001101001111110001010100001100011000010110011010000010101110100001010011000101100011100101110111010010011111000010001100000001001101111111011001100001110011010011110110100011111010000101100010111000100011110111110111100001110110100101100011010110111100110110010011010011100011101001000001011011110010001101101100101100110011111111100111010010101011110001101100001101100001000001101100101100001101111111110110001010010000000001100100110100111000100110010111011110001001011011001111110011000100010010110100010010101101101010110111100101000010011101011101100111000011011101111011101001000011001010011100011101100011011010100010110000001001101111101001110011001000111111101110101100110111000100100001100010010101101100110001001101000110010111101101000000110111101110111100110000111010111111111001111100001110111000101101010000111001111010000010111110011101111010010100110001010100010001001010011001010110011111111011010111101111110100101111111000111010101110000110100000101110011100111101101110111001101011110000100001000100100000011111011011101100111111010100001101010111000101001000000101111010011010101110100001101100110011100001111000000101001001111111101100011101001000111101111111001011011001101010011111000000111001010000111010111001010000101111101010110001111000001100110110110011011011101100110010000001111001111110000111100011011100111011111100100000001000111101000110110101010001111000101011110010101011000110010101111101000101001001110100100011010011001011110011010001000011001101111100011011010111100000000000111110110000001101000100001110111010100000010001010110011111100000101010111101110111001011000110101001011101111110010111011110000010000011000010011000110100101010010000010111111001111100101110000101001111001101100011010101100001110111101101100011100001101100011011110111011000011111101100110100100110000001100001101101011000011111001100001011101110110001111100011001100010101100100001101111100011111100100010100011001101000110100111010110001110000101100110101100010010110100100111111110111010000010001100011101001110111101111110100110100001010001010000000010100010101000010111011001111001000111100001001101101011001111111100000001111110010110110100101001001000111000011111111010100100111010110000010001010101011101110001010000011100010111001010111001000100000010111101110110110000000111010101001100000001100111011100011111111001101001000011100111000001100001110100001101110110001110111110001111000011011110001011011101101100010000011111101111111101101100111001101101100001001100100111110001010010100010011110100110011101111111101100010101110110011101010000001110100100011101100110011001100000001001011001010101110101101100000010100100011100101110111001111000011011111111001010000111001111011010011110100010011001110010000001111001111011101111011010100111111100101100111001100010001000100101110110111111011001001000101100010000101100111100111011101011101001000010110101110100110011010110101011100010101001010000110111011110001001100110001010001101110100000011011100001001101100110000111001101011100110111111110011110101010000110110110011010011010011110110100100001111000101111111101000100110010111101011011011101011110101101011000000000110001011001010010111010100001100101001010101000000010101011000010011110010010010101010000010011010101011011110110001110000000001111110110111101010100101110101101010001011000000100111111110101001010111010001000000000110010111011001001000111101110101000010110100000100010111110011000100011001010101100011010010110111000111000010110011110100100101010001011001111010101010011000111111110110011110001110001011110101010101001001101101101010111001100111010011110110110001001110110111010010010010101101111011101110011001011101011011000100011111000100010010101100000001110111101110010001110011111011101110010111110011110100110110110010101110010111001000111101010010010111000000101100010000110111100001001100001101001111011111100000111000011100100110010101001110011000111100011001010011100101001000000111010011011010100000001101000100100010110110010101101101001000110011011110000001110011001000110001011011110101111111110010100100011110110011100110111111011011111111111100100001101100011101011001001011010101110011100010101000101000100111100111110011111111110001010001001011000010111010101100001001011001010111010101101001001011001000101111110110111111110111001100101111011100110101010001001111111100001001010110101101011110011001011100111011001111011011001001010110110010010000101111110110110110000000010001100011011011110001101100101100101110010110010000110011111010001011111100011011011111011111001011101101010110110010110000101110001100010001111010100101011010111111111100100110111001010000011001111010000011001001101101000100101001011111001101000101100111011101010101110110010100011000101011001000010101011101110010000010111101100101010101011010111100000110010101111010011101100010011101100010101110101110010100101001001011010111101000010111011001100011110011100001111000000001100011000011100000001000111111001010000101100111001000110010010010111001101001101010101001011011110100011011001110010101100111010111011111010001001000111111101000001001100110011111010101001110010101110101000111110011011100001001000111111111100001100101100000100100100000110001100010000110000001110110000111101100010001011100101100000011000100000100101111111000101001011111100010101011001101111110100110111000000110101110011000100101110110011011001110100111001011111110001011001011000100001111010010111010111111110110101110011110001101101101101110010111000101000000100110001011001010000001111101000110001111001000011010010110010110000010010001011111000111110100100100111110001011110101111111100010101100111100110110001001010000110001100100111101111110101001010111101000110111011010101010001001000111011011001111001100010010100101110011111001101000011101001010010000100111101010000100010001100110100101001001000011110101010110000100111000010101010100010110011000100100011000000001110110010110111001010101111011100111111010100110110010101101010101111101101101101110110100011000100110100100100000011100000001001010111010000011000010000100011101100001110101110100111100111000111000111100110001001010111110100110011000100010011011000110111101111000110011010101000101000010011101000001100110011100100110110111101010100101100011010001101111100100011000010000101000010010110100001110011110101111111011100111100010010001110000111011101110111011111101001101001110101100101100110111110101010110011001001010111001000000101011000001010100010011110000011000101101001111000101001000011100001101111010111101101001111101111111010011001010110001010011111111011100101011001101011000011011000111110100011011011001001111011110100011101000001001110110111110100000011100000100111010000000100001010000001100100101101000010101111000000011000001110000101001111010111111111001001010001010001111010001111110011111100000110110011110011100100011111001000000001110101010111001000001011001001001100011001110010110111001010101000001000100011100111100110001001011011011100011011010101001110101001101110101010011001001010110101110110010010011001110000111010101100100110001010100011001110010100011001110110111011110111111010010011101000111011110110000010101000001011111101001010011111000111010010101010101100110111011111011101011011110000100111100000110000001000101001110010010110100011100100110000011000100001111111001001101111000100010010100100011011001000101001001111100101110011100110010101011111011110010101101010010001101000011000100010110100001111100010011000111001010000101101000110101010011011101110001000111110111010011110101101111000100001111010010100011100010100011111011001000110010101001101100001000011001011000011100100001010011001110001110110111010010110111100111010111001100001110101010011110010101010000101011100010011011100010101010011010011000101101011101101011111011001010110011110001010001111101011100110010101101101000001011111101010010101111110000111001100111111011111110010000011000100011111000000000010001110000010101001101110101111111010001101000011100000110110100011100100100110010010100110101001100101101101010010011110011011101001000111111011101100101010110011111101101110100010111000001110001110101011100100011011011001111101101010010101101001111000110001001011011110010000011111110011110111100000011011011110010111001001111011100000111010101000000110000101110010010011011010000010010110100001101101000001011110101001101100101100010001111100100001100001110010100110000110100100110100011100101011101110001101111011001100110101001100101101001000001001100111011111111000001010010011001100101100010001101111101100010111011110111001000000101001101000110110010111010101110100100000011011010001011110101010101011011110100011111101010000001000111110000111100010110000110100010001011001111110100000110011011001000100000000001001010100001010111011101000011010011111100011101110100101100111110001000111000011110100001010110011011001110011110100011011001101011110111000010111001100011011111111101011110111111000010101110111101010000010010011011000001010111010011001011101011000101100111101110110100101011000100110011001011001011010000001011000111110110111011110101010110011101111011111011010110011000110111100101011001101010001111110100000100101010000101110111001110110110110101011100000110011000110100110000110011001100001111111111100110001100011110000001010000001111001011111001101101100011011111100001001010111110011000001111100101000101000101010000000100100111110000101011101100010110100111010101101001100010001010011011101111001110100011010110101110010000010100110000111001000001110011111001110000001100101100000000001000111000011010011100101101111011111101111110110011110111001100100111001101111101110101001001010000101110011111110010010011100111110101011011001000111101001110101101010110010100000101101111100011100011100100000111001110100010000111011011000000001010110000110111110101000010100111100111110110001100110011100010110101111100101101000000000111000100111100100011101001101100001111110110100110001111111010100010111000000011010101010101101101101101000011110110101111101000001010010010110011000011000011101110100001000111001010000011101100010001010001001111100001101100001000100000101011101110110101110100011100000000110111010111110000000100010101110110001000111010100001111110110100000001100111111110101110010000001100110001100010000011001001000010110101100011110001111111110011100111000101011100101110111101111001001000011010011110101010101100100000010110011011001010101011100010000111000001111100110000101111010101110011001011100101000001001000011101100111000011101001011010100111001101100111011110001010011111111100101111010011001011101001001111001011110000011101000110111110000001000011001010101110010001011010111001100011111010101000011110100111101110101111100100011010111101001110110100000111000111110000101011010010101100110001000011100001101110101010010110000000100010000111101101111110101000101011101110101001101000010000110011111111100010100001011001100010111000101000010001110000111110011101001001000001000011010001000000100001110111001010110001000001100100100001010111010111001111001010010000111110101001101111010110100010011111100011000000110011110110001100100101111110111010111000100000011010010101100100010110000000100101001101111101010110101101111110010010010110101111000010100001000101010000101011110101110011110011011110100010011111100110110110101010100101101111110001101000011101110111110101111101011111000110101011101000110010001111011100001011010110011111001010010010101001000000111110111000010010001011010000101011010101001011101100101110111111011101000110001110001111010001001001011010101111010001100000111010110111100101111011011110010101101001001011010001001000011011111110011011100010110101000011010110010011011110001110001010101000110101101111101111110001101100101010001101111000011100101001011000011100101001111110000001101010011001110110001000111100111111000001000100000111110011010001100100101010000000001100111000001110100111111001000000000000010101000001100100001011001110110101100001010111100101110100100000011101001010110111010100110101101000101110100111111011010010101111111011001010100011101101110111010010100001000111101101110010011001000011011101010100011010011000111010000101100111111011011000101010010100100110011010011110110000010101111010001111001111001010010000000100001011000000000000100000110100010110100110101010010100111001101100001001111001111101010011110110000100001000001011100011100000110110010111111000000010011011100000111110110101101101011011001001100101111011010110011000110100010101100111001000111011011011001101101010100000111001010010001000010010001000101010000101101110000101011111011011011000011001110011110110101111001101110100001101110010000001110011111110011101001011000011111100100010010111110110000110110100110001001110001110000011000100110111101010111001011001100111100100111010100001010001010001111101101001001010011010100111111000110000000000100010101010010011111101100110101001111111011011100110111101000100101010100001001101110110111010111001011110011001001111011001011110111001100001001010100010110100000011100000001110100111111011111110011000001110010111010011001001111010011010110010010000001100100101111010011101011101010110011111100010101101110000000000100111110101000111111110001100100011110111001111101000010010010100100000010100001111011101011000001010011000000010100110100100010000010100100001101111001111011010100001010001000110100111110110110111100110101011100100011100100010010010001101111000110001101001011011001101011000111001011000001011000100000010010111110000110010110000100001011100111010001101111000001100111000101100100111101100110100000010110010111001010010101000001110001011010110110101111001101010111010110000000110110111001010101001001011011101010111100000110000101011000010100001000010111100110000010010101110000011111101111010000110011011111000000001111011011000010000000111010010110010011000011011101101100000001011011101011001011100001011111001101010011010110110110000110010101101100110010000000001101110100110010010111000100110010010010110101100001100010000100001000110100111011100011111000100011010000110101111010110100000101010100010010000110000001110010101111010011101100111001100011011010001001111011010011010010110100100101011100110000100000010001000010111101111001100000011000011101110000010101111000111100111000000100010001000010101011001001010111110001100010001010011001001000010001110100111111111010100011000110100011111110000101010000010010100010111011100111000000110011101010111110000010100010110110100011110111001010011010111011001101101100011111100001110001010100110100000100101110010101111111000011100100010100000001100001001100100000011001111111001000110001001101111111010001011000000111010110100110101011100001100011100111001101011101101101111111101110010011000101101111100101000001001110000001101111000011101100100111101110011011111000001100110101101110110110110011011001101100100010111110101110001110110111000010010111000001011110111011101111000010001110100111100101011111010110000100111100110110111101110011111011010001011100111011100100100100001100110101111111011101101111001100111100010011110010000011100110111010001011001000100110011101010111010101000011101101100111110110010000001011111110110010111101101111000001100100100110010110110100111111100100001010110000100110000101000101101011000011101111010000010100000101001100111001011100111101111101000001001100111001100111100011010011110110000110100100011100100011000010111111000100111110100100110101000110000001100101101101111000010001010100000101110110010110001110101111101111011101111111101010011011111001001000101010101000101011101101010100110101101101100110010110100001101010010110010000110001111110011001000101011010010110000101101111111010111000011111000100111111101001100100110000010110011011001010000101000100011011000100111011010100010000111100000001111001000101011001000011011010111010011000010100000111111000101110010111100101100101101010001111111011101010010010100001001011001001000010011010101111100001101111011000011100010101111100111001101000111011100001111111011011001101010000100011001100001111111101000101000101011001001010001111100011100000010110100111101010000110111000110101110100000101000011011110001101110111111000111010001111011111000110100010000011110110111010010111011011100111101111000011111101101000111011111011101100111101110101111000111001100000000110110111110110100110010111111001011110010001110110011110111000100001001101010000000100010000000111110110111000111000110101111011101100001001110000111111111010011000101100100001110011111110111101100010100001100000100101000011101001110000101101111101011011000010110110001110011011011000110111000100101000010010110110011010010111101100110000001010110111111101011001000010000011110101010010010111111010100110111010000111111001100011010010111000010001111101001001101001010001100110001011111001101101111010010111010110000110101100110101101111101000110011100011001101101101000001010000010111101111110101111100111011100000111011011101001000110011001100000111000110010001100000011101111011100011001011101011011100000000000100010110001010100000110010001101011000010111100101110110101011110111011000111001011111110010110001111000010001110101001001111111011011100111011000100100100110111111100001110001001010001101100110100001101111000011110100010011001111000110110011010100001001110011001010101000001100011101001001111111000011100001000001110000101011111011010011100101100101101101011110010001011010111000101101100101111000110000111111110100000110110001101011110111010000010111110110100001101011111011111011110001111011110101101001110000000001101111010100000000001101101101011100001010101111111011101001100011010000101011010110000100001111100100111111111000011000000010010001000011101100001111110110001001110110110000111101100000111101001101011010001011011010000110101100001100111001001101111000011011011001010100000010101111110100011111011110110000111010100001101100011101111001101011100110101111010000111100110100001110001000100010001010010010011001001011011101011000000110110110100100011111011110001100011011110110011010001001100001100001000001110001100000000100110100001001111001010100010001011000000010001110010011000101001110110011010011011101001010001010011001000000100100100100011001001111010110101011111001001101000000101011011000101110111001011111011100001000011111000110010110000001001011100000100101011100101000111101000110010011011011110010001110101100101011011111100110000011000011000111110111000111111010011000101011110000011100111010101000000101101000110001010011111000110101010111110010101011000010011111101010010010111010000000100010000010011010100011011100111101000011110100110100111111000100100001101001111101101100001000101011000001101001000111100010001111001000010001010101111010000001110001101101101010111001010001001001110001001000110100100100111000111111100100111000101101100100000010011111001010100100011111101100010101010110000001111101010101001101010110011100011000010000110110101100101100101101110110101101111000111000011101001110011110100001011111110100100010000010100100101010000110110110100010100001010111110011001001110100110011011010010011111110101110011000011101100001100001011001110011001111010110001010000010011000110000110110100011110110100011111110101011010010000101000111111011011011110110110001011110011110000001101010011100101010011100111111001010100101101001011100110101001010010000011011110110000100110001000101100001101010101011110111110100110000100101010111100000111000011100101110000111100011000100010101011011101111010101010001110000101001100010011011101111000101011000110001101111101011101110010110001001100001101111110000111000101110100001010110111001010111101111101111110100110111010000110110110000101010000001001011111001100111100010101011010011001110111011000101110000100111101101001100111110010011010011111110110100101110110001101100100001011000111110111010010000011001111110101000010001110110011011110110010101011000111101001001111011100101011010100110100000101111111110001010011100010010000110011011101101000101110110100001010000111100110110101100100111010111100011110101110011010011010011000100110011101001101101101010010000100100000110101010010001110000001111010110001011101110001010111010000101100100001111011101001101010000110100111000000110101000110101101100110011101011000011001101111000100100111011001110110011001100001000010001011001001101010011110000110101001100001110101110111000111110000100101010000110101110010011000101100111010110001100110110101111110001000010010010111100100000011001001011111001100011010010111011100010101100010110010111001001101011101111010101110001000111000000111111011110010101111100111001110110111001111011100001001010000100101001111011111100000111100010001010001001110110011111100011000101111010110010110011101010010000111000011110001000000101011111100111000110101111010101101000011010001010110111010100100101001011010110000111100010100111100101101101100100101111011011111110011111111110001111100111001011111100001110000100100101000011101110101110111111101000000110100010111001100011101000110010001111111100011010010110000101000010011011011110111101000001001001000110010111000001000101001010000100101010110111011111100101110110001001010101110111011110100001010101000101111001000000010100111001001010010111001100111010100101011100101011010100001101000100001100000111100001110011000011000001011111000100110100100111100100010000011101110001101011011010111100110110101001110111111010011011111100000101111111100110100011000100000001111110101110100111101111010100010111110111010110010011101011001011110001101100111000000101000001110100110100100100110110010100001111000010100010111111111111110011110010001011111000100011000011011010110101011001110000100000000011100010010011000100101110100111100011010010000010110111111011000000111011100001101111000011000100100100001110110010111100010110100111010100101001010001011100011110100011110110010111011110001000011000000010111010111110111000000101101001001011101111110000010110000011010101100100011110101011100110000000011101101000010110010111111101010101110100111111111111010000010100011000100111101101110001110101100010101110101110110011100100101010101101110111100000111010010011110101011000101001011100000000101010111111111100110001110011111001000001111000100010110101001110011011110111010000010010101011111110010000111000110111100010011111100111011100111110010000101110000111101001001111111101110111010111111101011101101101101000011101000011111101000010101101101101001110000111100111001001101000001000011101000011011100111110001011011000010100011110101010010100001110110111110000111110010110010000110110010000100100011101000110110010111101110000101000110110100100001011110011000011100000011110000000011100010011010101101101111110010110101111110110001010000110010110101010001101101000110111000010000110001100100101110110111000011101111110111111110111110000001011100110101011101000010100100011110110011111011101110101011010110011000111001100011110100010011001000000011111010010111110001100010100110011010010010110101100111110011001011001101011000111100100110000000111010000000111010100010111001111100100111001001011010010000111110101011011010101001011111110101001101010011101101110100010001101100000011000011011011001010101111001010100111000111001000001111101100100111111000010111000001000010111010011101001001011001010011110101011100111000001110110100101011010001011111011011111010010000111100111011110101110101001100001110100101010000110110111011101100000000100111011100000100001101000010000110111010110000101110011000101001111101100101010110111100101001010110101110101001001100011101001000000111101100000011001000010001011110010010111010100110110100101011001100011000011110101010110101111110101110001110000111010111111111000000011010000111011101001110101011010011100110001101101000111011001010111111011010010011000000000101111110010010101111110111000111100101000100000001010111100010110110010100101101010110011110110111011111111000110111001100110010010010000100111110000001110101100000110110001010011101110110111010101011111010111001110000011001001111010000001011011101101001000011110010011110010011000000110011101001110100010010110100000100011011000110100110001010011010010000000000010000011101000100100001011010011010011001110110001101001000101001100011111101101011110000110010011100010010010000001111001010011101101011010011100101000011100100100001100010011001100111100001001000111110001110001010100011100001100001101100000111111000000110100100110111100011111010101010100001000010101110010110000001101111010010100101001110101001110101000100100011001011011000100111101001000110000111010010001001001101010000010011001010011001100111011001100001111011100110110011101100110010101101011110101101000000010000001100010010101000010011000110010011010100011000111010000111011110101011010000100010100001101110101011001101001000100000011001011101000100010001101101001011100111100101111100111000001010001000110110100101000011101110010111011100111110001100001100100011110110001010101101100111111101101101000101110110110101011010111111110110101000101011001001010111001010100100001001011011011101111010000011100011001100100101000101011010111100111000100111101110101010101111011011111110111101001000100001101011110111100100011110100101110100100101000100000101101000100111010110110000000110011000111111111110011110101101100011001110010101001100001100100000011011001100001011111100110101010101000110011111001001110101111100110110011100111110000001010011001001100101000010101111011000111001101001100111101101110010001001101000101101101100000010011010001110100001100110000001010011001000001100011010101000101101101011000101101111100111001110110100010111111001100001110111101100101110011111101010011100110100111011110010101110010011001011011010011001100100100111010000100000110111110100011001011100111000101000010000100110110010101110100010001101010101101011001000011011110000011101010110011010001011011110100000010000010000001111101111100010101100101110010100111101011110100010000110110000001011101111100010011010100000011011000001100011101110111111000110100111100111001000001111000011110111001000100100111111010101001010110110110011111011001010000010111010101100100101001010011011101001000101101000010101110101010101101101010110001101011110101000011010001100011011111011111100101011101111001111000110111010001010000001000011011101011010010110110011011010010111101011111001010111011101000001011011110000011110010100101110111011101011000010000101100100000101110101001111101000100101001100010110110011110110001000001011000010101011001110101110011010111111010000011011010011101010100101100011001011101000010101000010101011001011011101101000011000101011001011110011011011010101110110000000011001101101111011101000001000111111000111111010001011000000100001111011000001111010111011101111001101000100110110100011010110000010111110001101010010011001111100100100111011010011101100011001100001011110111100000101111110001000101011010010010001001001100110101100010000010101010011010010011111000010101000110101011000011110001010000010001011010100111100011010101011111110001011110101110110000000101100001110011011001011110011110000101010010010010100101000101010100000111000110000010110011110000010011000000110010110011011100000110111010101111000100101101111001110010111100011100001101011000011111111010101010111111000010001100001000000011000100011100100101001110010010110000111101101011100001001101110100001011011101111011100110010111111011000100110111011001010111011000000110000000010011100011101101010100010101110100011010100011001010011000101000011010001110011001100010110000111111101001010010101110100110110011110101010100111011110110110111110110001010100110101100101100010111000011111101110110010000011100100111011100110001010001110101111110010011001011011101111101000011001010011000011010100000111000101101010001101111111111010001110110100011000001111100100110111110111101001101010100000010000100010111001110101101111011010110111110100100000011101011101100100110001001100001010000000011101000100100100111010101101101000001100100101010101110001111000000001001001001010100011101011110100000010111000011001110111111110100011101011100100100110000100111000110110011100000000100011010011010100101111101011110100001100110111101111011010111000101110111100011110000101111100000011000000000011101000011000011001101111111100011000101001100111110110010101000111101111111010011101011111101110000011000100111111100101010011011011011100000110111111100100111100111110100101100100111111000010100100111011000000110110000101001001100000110001101000000001010010111001011010111001110101011110010011111100011011110101011010101011001000110010000110100111000111100110011000010110001011100000111101010010011100111011011000100001110010110100101010111101010000011110100110000000111001101111001100111010011011100101101011111011010011011100000011010111001000001000001000110111111010101010111010001011010010011100010011000110101010001100111110110001110001111011010111011100011011110011110101001101110110111100100110001001101101010101001010101111100001000010110101100010010001100110010001001010001110110111010100100110110000101000011110111011100000000111111110101010011101101100101010110000010000110101110111001100110111100001010101101101111110010101010010010000011101000111010100011000010011010001110100011110110111011011010110000100010111000000101101000001001101000110100110000010010110100110011001100111010111000110110011001001001011001011110101100111111111001101000101011011111111111000001011111010011100101111001001100111110111111011001001010110010000011010101101010000010010010100111111100000010101000010100101011000001111110100110100101000001100110011010001111001001100101010011011000000011000010011010011101000100011101011111001010011001000111100000010100000101110111110001010011111010010110111001110110100010001100100101010001111001100111110000111000111010000100011111100001101110110101110000100010101010110000101000010111101100101111001111010111010011011001010101010110001001101110001111010000100001000111001001100011101000110000101010010110111100001110000001001011000110001011110010010011101111100010101001000101000011111111001011010000011001000101100101111111111010101010110010100011111100010000100110110011010011001001000001101110111000101110000010011011011111010101101000100010010010011100000000001010111000001010011001100010010110010110011010001001101000010000010011000100000001000111111101100001010010101110000010101011011001101000100101101001010011011100001011110000011101100000110010110111110111011001000011001111011011100110111010100100100101000000111101100101011011001111101001101111110101001100010111011111100000011011110110111011001001110100101111100110010101110010111011000010101001111000101010001100110101011011100110111010100011100000111010110000001111110011100010101010011011100010110001101001000110100000011010001001000100011101100110111110111101100000010110111110001100000110110110110000001101100110110011011000100100100101100001100011010010000000111100100000000110001010000101110110010011001010010110010001111101010100000000011100110000000100001011010101100001001100110011001011110110011011111111110010011110000111010100010101101100101011010101101110101010110111111110110110000110000001011011010100010101100111010110101001110101000010001011110101010001011111000011001000111100100110010000110110000111100110110011000010111000010000000010010010001111111101110010000010010000100000001010010111001100000100011001111110001001000110000100100100111100111100010100010001010000001111101011111111100111001111010101110111111100001111110000011110011110010000110111111110100010100010010001001110101111010000111110101010000110001010110100100111110011001110011101111001110000101111011011000111000111111011111100110001000001111111101111111011010000010010111011101111001101000010001000100101111011010010100101010101110110110110011111100111001100000010101001011001000001110110101100110010011100111101111000100001100101100110100111111000101000001100110110011010011010000000110100101100111001000111010011000101000000011111111011011011010010111101000000110110001000111010010101011101101000000011110100111001011010100100110010100001100000110001000001011111010011111101001100010001101110010011010101000011010011000001110001000101000000011010011110010111100110001000100000001011010011111111100000010001111100100000000011101110011110000100111110001100101110011111100000000110001001001001001100110000001100011100001010010100100110101011011000001001100011110000001001001001101000010011100000001111011011101101011000101000100000010101010111100110110011001010000101110100110000011000110101000001010101011010111101010100000111110000111101101111100100100110101010000000001100111010010001111000100110001011111110001110101000010001010111000111001001100011011010100100100111001011011000100111001110101010100110111110101110010000101000101010101111111001101000110011001000011001010010101011110110111000010011011110010111001000101110011100011110111101001111011100001010100110111010100111111010110011101010100100001000010011111111110100101000001010110101000010010100011100010000000001001011101101000100110110001001110111110100010010011010001010111111100010001110100111010001110111111101100011100101001110000100000010111100000001110010011101111111010001001111110010001000010101101111000011001111101101011111100010011100010100000100011001111111100010101000101001001010001111111001001010110001111110011011011011011010011110110001010000011011000010100000111101010010001011100100010011111110011011011000111001000101101101101100111001111001001101111001110100011100101111101110111000010011100000101101001110110011011000101110010111011101010011000000110100001100110101100000100101101000010000011000010110000011100111011111011100011100011111011001000101000001101101001000000100010010001101100110101110100000100000110010100110110011110100100001100111000000000101000001011000101011000010001111101111000000001110110111000011010011011111010001111010010011111000011000110000101111000001111101110111000001001101011011010001010011011101100011101010011000011011100111111100010000110000111100101010000010111010000011101100111110011010000011111111011010110001001111011110100111000111101110011101001111110000000000111000011101111100110010011011000111111000100010010000101011101011001010100101100000100000011111000111111011000110101011010000101101010111110110110001000100110001011000100000100111100011101100000100000001110001100011011100011010000010100010111011111010111001000000010101000001111010011101110111110010010001111011010111000101100011011101010001010011011011011011100110000001011011011100001110011011001111101011100011101000110111101101101111101101010111110111100110111100000001011110010100000000010000001110101111111001110111010100011010100010001001100000110000001011010110001010011001010111001100110011001111011101011101111100010001000111011101001100111001010100111010100111100111010101000110101101000011110000011110100000010001011000110100101010010001101011000011110110110111001010000110100101101010110010011011111100101101111011001101000010011010110111010000011101010011101110110111100001001110101011111010101100110010110110010110100001000101111000001011011000110000101011101010110001010110001100110001001101101111001110110001111010110011010100100100011000000110110100101001000001110011010101100001011100111011101111100110011100110111010010001100001100111001101001100101111011101111001010101010111111010111101111011000101001100111010111100011001111010010010100010001000100010010011100111100100001010111000100111001111010100110111111111111111011110111100001011100110000100000100111111111111111001100111001111111101110101000100111011000100001000100010010111001100010100011000010010100101011110011100101100101110111000010000101111101110100110111110010011111110101111000101101011001010011010100110010100101011000111100000000100000010001111100111011000000011000010010110001101111010101010011011100110000001111011101110101001101101011010110000100010000000010101011101100101101100101001100011101000011001000110110110101100001011111110001000110011011001111101111000100011010011101011001001010010010011011001110101101111110000001110010010111110010101100010001100011100000001000111111110101001110110101110101000011100001000101110000110110011011010100000110000011011000101100001100111000101100111110000101100000001011111010001000010001110101001101101000111100001011011011000111100000100100100100111111000010111110011011001110010010011001001101100101010100000111001111111011010100110001111110110110111110000110011100010110110111011101111111111100001011101000011000011000110010100110001010111110001111011001111100111100011110010101011001100011010100101001100101111110011101001110011111000011111100000001000001110000111011011010101001011001100111011111111110110110010011000010001110000011011000100111100001110010010111010010000010100101101011101010110001101110111011011011000100011111000010001011111110010000101010101011101100001001011101100101111111111010110001010000110000110101100001000010010011101000110100010111101110110000100111101000101011000010111010111000110101010111011011001010001101110010100101000011100111001001000011110111010111101100101001100010101100011100011010011001101000000100110010111101111111111110100001100010011110000100011110111111101000110001011101100011010101001011001011100101010011011100011010000101000110010110111111010000000011101000010110101111010101110110010111010010011010011101000110000011010101100101100001010011010110111010011001100000111000100101111011101111111110111011111011101000101001010000111011001010010100100111100011010011011000100101101001101011111100111011100111001111111010110100010000100110010001010011100010011111011111000010110110011010111110010011100110101011100110101000111000100110000111000110011011111011011100101011110101101010100010010100101001100110011110101110011111010001000011101101111000101101000010000011001011011010010100110111100100001100100010000000001001000110111011000110101110011011001010001000010000001001101100111110000101000011100101000001111111000111100101101011011000011011101100010110110010110101010001010101011010100001101010010101001011111000011100000011100000000010100101000101101011001111010101100011111100111101101001010001011100101001101010010101110111110110010000000100000011100101110110011011010101100011110001110011000101101000011101001000110001011111100011100011010101111010110000101111111010101100110011110010010111110100110010001110000001010000011011010000101010001110000010100001011010011010111100000110101001110111010000101000010111011000010000000010000110010000110001101110101100011111110011110110101111110110000011101000000000001001010000100000000110001111100001111010000001010101011011110101010010100110010010111100011111011101110101111111101001101011100001001001101100110001111001011010000001100001000101101111110111101010011000100010011110110011100000011100001111001101110101000101001100000100010001111010011011110000000101111110110010110010110100000010101010001101110100111000000100110001011000110001100101111110111110011001101001100100100100110111001001010101010000101000011100100000111111010011100001111011101111100111101001111110110100100010100110110010001011000111101101101011110001000110110011001001011001100000111100010001101001001110110011111001100111000001001010000000011101000110010100011110000100010001110111010000111001100100101000000110011011001010110110001001111000000110011000000110110101100110011111000010011111101110010000101101001111100000100011111001100000111100001101010111101010100100001000011100111010101010110010111000101010010001111000001001111011010011001010101000010011011110110100001101001100101110110010001000010110101111001110101100110101001100100101101101110111111001001001110110111011010101100100101001111001101001000011001001111000011000011111000010001100101110001011011011000000000010000010011000010111110100111010000010010000000110010010111000111001100011010000111001010000111110111111111101100001100110010111100101111001001101001010010001010011111001001011101011011111000000101001010110001000111010110101101011000011111010000111001001110001111010001001011101100011110011101111010111000011110111100000001110001110111010011111111010001101001111111110111001111101001100111101001111010101111111110010110000011111100010111001010011001010100001101100010101010001110100100011101110111111101011000011111011111011110001100011101110011111111001111010000010000011011000001001110111001111101001001010101101001111011000001110101010011100001111000001010010000001111111101111000101010010011000000000100110011011001110000011111111101010100001011000111000010001010100010111100010011011111111001010000010111010001000001000011111111010000111111110110101000101010000001110101110101001101101110011010010111100010101110100010111000011001110100110110111101101110001100100010111001011111100011100101100010111000010110010001001011000011110010100010100000100101011100000010100000110010111110111000100010101011101111010001001101001000111111011010110100101001000001000000111110010011011011100001001000011011010100110000110011111011111101111011001101000010011001111101101000010100000011111000110110111001000011001000001100101011110100010010000011100011010100101011011101100101111011000011101011000110001111100010111101111001001110011111110100111010011110011110011000101010010000000001010100001110011001010110011011101111111111001001101001100101000001111110011010011010100001111110100011001111100001010101100001110101100100001101100110110100011011010001010001100011111011000100100011100110011011011100000101010000101001000100101001000001100000100010110010010010111100011011001110001110001110101111110000011110111001101100011101110010000100101011100000011011101011010000010001100000100101101000010011100111110101110000100101000100100101000000111101101100101000111010100111011001100110000100110100110011110110101111010111011011111010011100011110110101111010010001111110000101100100111110100111001111011100011101100000000100000000011011101010000110100000100101110011100010000010101010110101010011010101111101000110110110100100111101011110011101101110000111100100001011010101010101000101101111000001110010010110101011001101011100011101100000000111010110100000101001011010011110100011110011101011001000100101011111010101111011111000100110101111110000000110100011011101000110001011011011010111011110000011111111111101001001000101001111100100010010011011001101110100010110111111001110101011000111010000001010101011011000010011111101011100011111110101010010100110110001011010101111110000001101101000100110111011001011100010000001001010000001000110111001110111001011101011110100000001001101011010011100010010110001001111110110000110111011100000111100100000011101001111001100110100110001111011101110101100011111110000011111001100010101010001001010010111100110011101111000110101010000110100011100100000010111111000100011111101001001101110111101001101110101001011111111010000111101010011101110000110101000011100101100100100000111110101011101110010001011000111001110000111101010101110010010010110111101000111110000000100001110000011111100011100100110001011000000110001110110001000101111010111100100010100000110101111101000101001111100111110011011101110001001100101011111001111110110111001000010011010111000011001001100000111100010001111010011100000101001010000110110011011001110010100100100110110110011010011101011011010011110010111011111111111100111011110011001111000010101010000100011100011011010011010110011111100101100011000110110011110001101100000101101111010110001110100101011100011101100101101011000111111001011111101011110111101001001010000111011101011000111010111111011001001001111101011111010101010111000111111100000010000100010100011000011110100101100100010100100100011100110110001010111111110001100110110101100100000101011000010110110000000010001000110110110111101011101100001001110111000000010110011001101011010100110000111110100111100001110100101001110011000010010001100111010100111100100001100100010111001011001011001011100110110011111101100010001011010100110001010100110001011110010000101111100101110100011001001010000110111101111001010110110101101101110101100001101011001111001010111011100000010111101001010100111100010101001000001000101001000110111100011111011101111100010100001100101000011001001011011110110000010001100000100000001111100011100100110110000001010001110100110001100001000101001010110100101000110111001000010110000001100001011001001100000100000101110101111111110011010011100000001100001001111011110001001101011100101111000101110100100110010001100001000111111011000000111110011110101101011000010100001001110101100001000110101100010100101111101101000001001001111011011010000101001111111011100010111000100001101011011000100010010101101111101100000011001100010111101010010111100111001011110000100011011001010111101000001001100010011011100110111001011001001011110110111111010100111011010110001010100011101111111011011000011100011010001110011011000101000101010000011011101100010100010110010001011110001001101100101010000000110001111110000010110011100111000011111000110001010001111100111010000000100011110101000111111001111000011101000100001011111010100011001011101000011100000101001000011111001101001110110110000100111010110101111101101001101110010010100101010000001000110110001101100101001101100111010010110101101001101101000110100011011101001010100000101101011111010110111000011001100010100001101101000000010100100111100000001101010010111100011000010111110111100011100001011011011011111111001111100110101110011011010000011111100100011010000110101101111000110000111100011100110110010010010000011000110110000101110010111011100001110110100101100010000011000110010101110111110100000001110101001101011110010111000011001010011111101110000011110011011011110110100011101101101001110001101001100110111010000010111011001011101010100100000101101010100001101000100011011101101111100011110111001101010100111101111110000001101111101001110111110101011100010001000101111001100001000000010111101000011010001000000100101011101101110100101110011011111011110101111111001011011100111001000110011100011010011011100111100100101000010111101010110011111010000010101110111100100001101100111011101110100001110010110101000000010101000111101100111001101010001111100011111001100110111010101010111011111110010011111111011000001110011001010010000101101111100110101101111110011010000001000000100110101100011011110001011100110101100000100111000101001001110101111101101101111111110011111010011001111001100000111110011111000010010011100011011110010110101011011101001010001101010100000010110001101001111010101110010011111000110011111110011101000111110100100111001000110100100011100011111010001100001101101010110101001011110111100010100010010101111000101011000110101000111111111101011110101001010101100011010101000001111000101101010010111001110100000000111101011010111101001010001111101000000111011111110100111000110111010010001011101110111110010110101111100101100111100110001100010000101111101001110111111000000101001011000101011001100011011101010100001110111001001011010101101111110111001110101011111001101100011100010010101011010111100010100111100001010100110111101110100110101010001110011111111001000110100100110111111111000111101010111011111011010001010100101011101111101100111000110101001000010010101000000101110110011110001001100110001111111100010010010000110011010010101011000110101001000100110100010111010011010110001100010011011000010100100010000000011101001010110010000111000110111001111100100100100001001001010101101010110001111001001000101011011000000101011001110111000111100000000111010101101110110110011110000000100111011000010101010011011011011110100111101001010111011001111000000100011111101001110000100111000001011100101010001100011010010100110000001100011100110011000000000001011011110000100010001110111001001010010011111001010001111110101001011111111101000011011100010001001111010010100010101101110000000000100011001101111010000000111010000111110100100110111011011010010110000000011110110010111110011010000000100111110011011101001001101010110000001111001100011001001101100100101011000100011001100001011010011010100111001100001100000010101010000011000010011010111011101100001101000100011000011011101000100000010111110111111000000011011111101010011100100010001111110000010111010000101010100101111001000100000010001111110100101011001011001110011000101001001101011001010000001001011001001001100011100010100100011000101011000110100101101001011111101010110000010001011001010110001110111110001100110010101000111100000000000011110010000000110100010110000110001011100100111010111110111100100000000011010011100101011000000010111110111001110111001111001001110010001101100010111011101000000111110010001100010100111101111101111111110010110100001000101010001111111111011000110101010111100110000010111010111110011000010010110110010101010111010100100001101000100010111100110110101111011111101001010100111001001101010101100000101001001110100001010111000110100010011011010111010001010111111010111110101001101010100100100000011010101111100100001100001110001101100001001100010111010101011001011100001010101110111111100000010000110011011100001000011011110011000110000000110110001010100100110100110111111000010111110101001100101010101111110000111011001000110010011100110001001001100000010111110111100001100000011011011011101010001100110111000101100011010011011100101111110010110100010110101011110000011100001011011000010101011100010110111011111001110000110100110111001101101010010111111001101001000101100011011101000101100010111010010101110111100100001001101000110010100010110001111011000110010111011111111010101111111100011011000000110100110101110011001001011000111101100011010010110011111011001001100101010100100110000001011101000001100010011100011010000110000011111110011001110101101000101011001011110010001011011011010101010111101000011111011110001100001101001010010011111000110001001101011110100011101101100011111111010110011111011110001010010001100000001110101110100011100101011011111100100101101100001001110010010111110011100100000110001110001001001010111001100011010001001010010111001010100011110010100000000100111001100111001111101101111100001001010011101011111111100000010010100101010011100101100101000111101101101110111101010110010110010110001100101111110011100110111111011101011100110100001010000100100101001111110010010001011011011110001101101010001101001111001100100101011110101101000100101111111111010111100001000100101011010001001001000100011101101001101100010110010110001101000000001110111100010110011000101011101000111010010011111110010100001001101011010111111101001100111011111101110100010000011111100100111011111011001101101111111110100001010011111010010111001010111001000011001000010100011101111101100001101001110001100001110010001111110101011010011010100011000100000101101100001001100101010111000110110101001101111010101011111010000101000100110101100100010101110100101001010100110001001000111001001011010111001110101000110110111110101101101110000110001011111011101111110101100011010111101000111000010000000100100110001101101011011100111000111010110000101000101001000011011000010100010001001011000110011100111010100011011010010011000100100111011110110111000111010101101100010011001111000001000011100011011100100000001100000100100010100111000010011101100000000011010111011111111000111110011001010100111000010101001001010011011110010001111011000111100011011011001110100101110011001000111011001111100110000100100101101111101011001100111111000100101010100100010100001011100000001100101000111010101011000011110001111010101110111001011011001010011011011010100101101000011100011111101111101101110001111001001011110010100101000110100110011110111110001110101000011001011101010110001101010000000111000001000111001001001001110110110010010101010100001000011001001010100001110111001111111111101001010010010001000011000110010111111111100111111011110001110011111111011101011000011100011000111011110011000111111111101001001011101011011011000111101011101001010000110010011000111010111010011011111110101101000001011110010110110011101100100111011100000110011011111111111000011100000100010100000111010110111101000110000111100011001111010011000000101111101001101110110101110001101100011000110010011111010000010100101100001110100001101000011001101000011100111101111110000101000101100000111100100000001110000011010100101100101110001000001010101100111001011001101110010110101100111010010101000110111100100001101101110100111100011000100101100001101001000011110101110000010001011111001011110001010000010010000110110111011000111011001100101110011111101010111001001111011100101100001100100100110011001001011100110110101100000100000010100101000001110001101000011010111010001111000010010110011101000100001010010100101101001101011110101000010110001100100101111100011000111000001110111101011101110100010011001100110010110111110101101110000111110100001110011000111111110000000001100011110110010101010001000111101000101000001111010000010100010011010001100010001111011100111011100000100011110011000101000010011101100110011111010110010111000011100101100110011011011010000000111011100010111101100000111100010011011110010101010100010010010010110010001001101100010110100000110101011110011111011110100110111111101010001100011011001110011000010101001100100011111101100011010010110000100001101000010000110101011100100001111001011100110101110011001010010000110111001011010100101101111010101010001011111110110111010010101100011000101011101000011101110101000110110011010110001110110100000011110101110111111001111110000010111000101110101000100000101111011111111111011111111000001000101101011110110011010101111000011010010000001000010010001011101100101101011101001100001101000101001111001110101100111110101001001100000010001011111010110111000011111011001010110100101011000110101010110011101100111000001000100111111110101110001100100110100010000101011100000001111011110010101101010100101101000001010001011111010000110010011101110111010001111000011001000110110011101110111011010110111000001100011000011000011001011111001100001110010100011110101111001011100000110011011111110011000100000100100001011110011101101101001100111001001111001111101100111110110001111111100100011111111000011110010100010101110110001000000110100110011000010011101101011011101110111101010011101101000000000110101010110110100110111100100100111010010010101110111101011001010100001000101011000100001101001111000011111100110011111111110101100011001001100100111010100011011000100101101010100010011110011011001010110011001110011001011000111011111000101001000000100011100111000010010111100011000000000100100101100110110101000110110111100100110101111100101100001001000010011100111100000100111100010010101110011101110101100100101100101110100101000111101111101011101111110101101011100111010011011101110110110010101011101011010101110001111110000001000000100011010010010011010001110111101111101100010101011100111010111000111010100011110010010011010011100011010000110001101001010100000000001001101000001100001101101000100111100011000111101000001111001011100011001001001110000010101101110101110011101111100010100001001100111110111100010000011111001010000010001110101000111000000011011010111111101101100000111100010001000100011011011101000101001100000110101011111101100001101000101000011110100000010011001011001011010101001110111000110101111010100100111111000111111010011101101110001001111000110001100101110011000001110101011111111000011111100101111010000001110100110100110101010010010000100011001011100001010001010101000110011101001011011001111100110110101111100000101111001111110011100011000111101010111000000110010011101110111110011011101010000001010101111001100010001001110111100001110111001101101110000110111011000011011000101010000001100100101010010000111101000111100101000000110001100111011111110111111110000000111111000001011000010111000111011111000101010100111010001101000101000001011001111100100100001100100101010100100101010100101011110111010111000110011111001010100000001010011100010011010101010001101111101001001100111011110011101100110111100100011010010110011000101110011111111000100100011111100111010001111101011100100110111011110000101111011110000110100110100100101100000110010001101111100011110110010010110111100110110111011111001011011010100000100001110010110111111110111100110010101000001010011010001010110100000100110100110101001011011001100101000110000011010011110101111101010101100111000101111111110011111101111111100100011100100110010110000000010011011110000011110110011110010000011110101010011100010111100101001111000000011010011000101111110011011100001100111001111111001010010101110001100111101011011110101100000010001111000110110011000000101111101010100010101101001110101010010010001001110010111101110001001100000110011101110000001110010110100001010101110001011001011011110000100001100111110101001100001010000000011110011100101000010011011011111101001001011101001011011110011100010000101001001111100001100001111011000100101001010111101100011010111010011101101111110011010110001101110001101011001000100111011001011101000011110100001010110000011100000010010000100010000110010010010101110110011011101111101000110010010010100001100000110010111011011001001011001010101000111000010001011101001111100001000000010101100100010001100111010111011110011100000010101010100000101111111001000101001110100001001011111001011011001000110000001100010100101011010001010000010011001000111110110011100000011100111100101011001000000010101011110110001110110011110011001101010101011011101011101101111001101010010101001100101001010101011010111000011011000101001111000101011101110001111110111110011110111001101110010001001001001001100011000010111101101010101000110101100000110100111101101101111110100000111000111000000110100110000011110111001010101001010010000011011010111101010000101010001111110110001001100101101001100101001111010110011110011111101011111011000101111011100000011011101010111010011100101110101000001011000111010001001111001000010101010011001110010011001100011001100001001000010000001101101000101111101000001111110011111110011110101101000100100010111011110101010001001000011000101100001100101101001010110101001100001111111110011110010001110011000110001110111100000010111101011101000101101101100110011011110011110001111110001011100100110101001101011001100101110011001011101010101110001110111101100001101101111110111100000111111111010001111010010001000111011011001111101101101001110111111011110111101010010010000101001010000011010100011110110001000100111110001010110010101011010100010000100100011001110011110001100010111011101100011101000001110010011110001011111111100000010011001110111010111001001011100100101111001100010100110101100001000010011111110110110111000011011100001011001110000100100010111110110100010010111100000110000001111011001010100100000010011001101001011110001111111100101001110100101110111010111111000001100111111010011010110110010111111100100111011110000010101011000111010100110010111101001101010101101100111111010001111001000000011111010011011101100011011000010110011101000101100101100010010111100111010101011000111110100111110010110111001110100000010101100110011000000111010101000111011100110000101000110000010010000110110100000111011010000000010001011000011011000010110011111011111000010011000100000001100011011100001101001001010110111101100000001100000001001100100000010000101000001111001101110001111101001000001001010001100100110001001101001111011100100111110000001101010010000000100111010001011011010110011101100011110001110111001001110011011011111110100011000111110110101110110111101100001100111011001001111110010111100110010010001101000000011000001101010001100001111100110000101100111011001000110001111010000101101110101010000001111001001111000101100010011000000000001100001101000111110110111110000100100001100011100101000100111000111001011010001001101101001001101110110011110111001100001101101111001110010101101011111001011000000110001001010101111000010000010000110011001111010000100100001111111010001001110110101101010101100000011000111000100000111101101111011101110010011110101001010011011011010101111101100010010111011100111110001010010110101100111100101011010010011000011111001000110101001100101001011101110000011110101100000101010101010001111011010000110000000000110010100000010110001010101101101010010001000111111110011010100000010110110110001010010001100101000100111001000100111000010100110100101011011111011111011011011001110001011111010000011101111101100000011010011110000100000010001010011010011001011110011001001001100010010100011111110000010101011111100000110001101111001100100000011011110011100100101010000110101001100000111011101110100010011000110111100001111010100110000000110010001000110111011111000111100100001010101101101100111111010100100000011010011111011100110110111101010111011010010101001010100101100010011100010000001111110001000110101100000111101011001000101111111101011111100100101011011010100101101011111110011111101011100010101100111001000111100100100000001011101100011010011000010100010101000100000000110001000100101110101100011010001011011111110001110000101011111011101000111000101100000011110111010111000110011011111101111110110100011111110011100001000010011110001110100001001110110101011010111100100110101100011110010100110101001011100001010001010110111100011111111001111111100000001101010111100010101111101110000111000011100000011100010110110111100110111001110111000100101001101000100100001110110010001110100100111010010001110001000011110010011001101101000110000110111010101110101001010101001110000111110100001000111000010111011100101010011011000100111110000011011111010100001000100011111000101110100110010010001101110011111010001010000000001101110101110101111111000011101010000010011111001001010011100010011110000110111000000110001001101110011011101000010101000100011110001000010111101000101010011011000001010010100000010011001101111110100100001010101111000101010010100110010010101001010011010000100000110101001111100100111011011100110010100110011001011111010101110101010111010111100110010000001001001100010110101011011101111110101110100110011111000111011011110001000010101011010011111110000010101111100010101111101011011000011110111011110000110100011001001010001100100110001000110011111101010000000111100011010110100001001001101000011011001111000000111001111100011100100000100100000101000111101010101100000101010001000010001100111101011001010011101010001011110000110001000011101110000101100000010010110011000100111101110110100111111110101010101110111000111110010010100100001111000101100111111111100001010011011001110100011110001000111101101111010000101110011000101011100111100011001111010110111101111111000000011111010000011100000010001001011011010010101010101001010010000010101011100101100100110101001000010100100111101011001110000101111101000011100100010101100011100110001011110110110010110011001010101101011010011000000000101111000101100000110101000011010001000101100001101110010101100101110110001101011111001111101011100110011001000110110010101110111010000110001111001111111010011010011011100001001011100111001110101011100001010001010111110100100000110101110000111001111110100110010110100110001110010001110011010000000011110000111001011110001101011010010010000110100100001011001011011010011001110000101001111011011001111110110100011001100011111100110110101011011011110111011111110111100100011100011010100111001000010110101011101110101001011011101100100111000111011101101111011001011110001110110110000111010111011110010101110010011110001001111010011110010011100111001000110100000100101100001011001111000011110001111001011111010011000101111100000111100111010101101100100101001110001010011101111000101111101101001110011101011010010001011010001001000110000100110011110010011001100001100001101001000011011101001100101110101000101110111111110100011110101100001001001111011101010101111010001101111001110101010000001101001110010011010101101100000111011111101010110101010001001011111001010100100001110101001111110011100111010100101010110101011111111111111101010000101110001000111011001001100111010010011101111000101001010010010010010001000000011101001111000110110010000100111010110010010111101000000000110100000010010011010000011010100101110111001100001110110010001111001101111111110010000010000110101111001101011101011000010001011110010010100010110000100001101110010110100011011000110111110011110111101100001011100101001001011100001000100001011111001010010110110111100001001100000011111111101110011100010011010101010101100010000001010101101110100001011000111000001111010110101000110110101111111011101001101111011110011011001100011001111100111011011100111110111110111111010101011111001010010110010010101010000000011110011100010010101101101000000100000111011100000100000001111000110011101001100101110000010101101001010101010110000101011001011001111110001100010111110001001110010110011101000001111111011000100101000101110110001110101110111001011001111000111111110101010100110100110100010101110010101011010010111111110001000011001001010101110101000100010110001000110001100100100000001000011101100000100111111101010111001110111100100011111011110101011100100001010110111011011010000000111011111000111101111110101100101000100001000011000010011110110000100101111010110011111011011010101101101110100000100000111101000101100011111000001010001011000001100010111001101000010100111110010100111111100001001000101100011101011101011100000110100101001101000110111010001001001010111101110110000100101011110010011001111010001010011001101000100000001111101010010101101111011010100010010000101100010000101011001100011111001000010010110001010000000110100011100000110100000110111010010110100000111111100100001100011011100001010000101101000001111111111000010001111110010001101110011101101110100100011100010111010011110100011100111100001011101100010010010111100100000100001001111101010001011000000111011011011000111011011111010010000111001010111111111110100101010111011010000011111000111011111100110001111111100011110011111001100010011011001001000101010010110011111001010100000100101101101111000000101111110001101111100001001111011110000000101011111111101010000101100000000000011101011010110000111111101100100111110011011001001011111011011100111011010000100001111000001010000000110000001100111000101001000111110101011100101101100100000111011001010100100101111001001110110000111010011010010100010011100111101100100111101001001010010010111101010000110111011010000110110000000100000110011101100011110100101110111010001111100011001001000101000010010101000111011100101111100000110001011111001100101101101010110000010000001001111101110100110111101101110100101000001011101011011000101001111100101100101110101010010000001100001111101111110101101100000111111110000100001111001101110000110110111011110101001110100011001100001101101001000011011110110101111110100011100000000100001111011100111110000001001001000000101110001010001111110001011111110011011010111000110001011000010010001110111101011100101100001110001011101110110010111101100111111001101110010010101000010101010001011110110101110010010101111000110100001101110011100110111011100110010000001111111010010010100000100111010011111011011101110111101111000001011101111000110110011101110000101000111000001011111100000011010000000111110011100111111000001100001010010111111111111100111111010100101011011111010011000001000001000011001001100111010100101011010111101110110101111111011000110000001101101011111001011111011101111011000101010000111001101111100011111001011110101011111010111000011000111111110111001011111001011000111100000010000101011110001100000101000000001100100001101101110101101011101101000001010100100000110111001000100111010100110011000100011001010001010110011100001000000111111101001010101000011000111010111111110110110011000011000101000010111101011001001011001111011110100000001110011101111000100000001111011101111110000011000001011100011010101100100111001100101101011010001111011110011100101001100111101100011010111100101011101101001101101100111010011110111111110100010001101010101100111000010001000000011001011010111110110000100011110010111111011011011001101111111010101110000110010110110001010111110010001011100100011010011111101101110100110001011111000010111110100000000010110100011001100111010100001000001101101010100000000011111011101111001010111011010110100000110101110101001100000001001111110111001100011011101101000110010111100010110010111110101011100000010110110111110001011101011100001110000010010101010011100111010100010000110100110000010011010110000111100111110001001011011111111100100011011111001100110011100001000110000111100001011010010111111011100110101110010011011100111100001101111101101010010011001100111111101011111000100111101010000110001000111000111111100100010101000101110100110100110110110101110100000001010000001000100000101000000111101010111111111100011101111010011000011010001111011000010110100001111000101110011000110110001001000101000010010011001011010110000101100111111110011000001100000100101101010000111100111100010000000100001101000101110110100011111001110001100101110010010000111100110000000100010111011100001100011011010111101000000010100001000101101001100101000101010100001100001100001110111000101111010100000011000010111000011110110000011111111000110000110100101111110111111001110011000111011011001100000000000000101101011110110001000110110100001110011000010100001000101011100101010000001011111010001111110110011001011011001001000000101001001001100111010110001101110110001110110100011010011010011100110111000110010001110111011101111011101110011010001101101000000000001100110000101100100101000111100111000000100010000010111011101111011011011010100111100101111110101000110010011001011000010101101001011111001100110000101000110111111110110110001111011000001101001001000111011001010010011111011011110111001101110001011111101011001110011110100011000101011011110011000111111010100001101010000110111011101100000110011001011111111001110000100010101111100000110001000101111110010001011110010110010010000001110101010001010100100010110111101100111010000100100000111010111100110110001110101110111011101110110001110100110100000110010001100111001011011001110101100010100111111011001010001100101011111010111100000110010101001111001101101110100011011011101100100101111000101100000110000100010001100111101110101001101111110110100111010110111101111001110100001011001011111100101011101110110101011101011000110111000110010010110011101100001011011111110101001101011001001000010101001011010001111100000010111101011001110000111111111111110011001011000011000011010100100010010101100100011110110110000100010011001011000000000000101101110100000110101010000001011011000110011010110101000101110110000110111101000111111101110010101010001001000101101110100100010100100110111111000001101101100010011100000110101010000011110010101011111010111010110001000010101010011010001010100100011111011001000001011110010111000010101011010011010010101000010010010101011001111101010111110100100011000010010110100001001000110011101011111010001110110000011011111100001000100111111011000100110100010001000000110110001011111011010110000000100110001100111001011011011100101111011010101110001011101100101001100011110001110001010000101101010100001001000010010010110110001111001110011000011001010011001011101011111111001011010010111001011011010111001100000111110110110111110101011111010101010010110110110011011001101111110110010100100010001111110100001111100010111111110011111110010101100001111100001110100011100101101010010110010100000110101001100001110010110011000111101000101110000101101100011001011011110101110100010011010110101010100100001101001000010010110111000110111011100001100001111100001110111111010000110101010110011100101111111001011100111000101110000101010100001011001101001000100000110111011110001011001011000100111001100000100111010001101011110111111111110010100100101110111111010011110010110001101110000010010001010101110010100101001010100001011101001110001011111010100000110001000000011010011100010110101011011000010110010110011010111000100110000100011011001011111110111111000000110101100001110101011010011000110011000001111110000100100100010101001101101101101000101000100110111010000011100110101011110110010110001101001110100101101001011100110010111111111100001010011101110011110110100000110111000010001111010110101010001111111110110111001101100101000101011010100000110010110110110100111011011100000110011100011010001000101100010100011101111101001010111001111101110011100010010100000010111011100001001011111010110100110101001110010111010001110110111010101100011100110100100010010101111011010001011001001101110010011010111010110100110011100001111000101001110101100101101100101010010001101000100111111110111010001010000000101000111010101011101011101000111010111100011001100100010000010000010000010000111111100101101100111000111001101000111001011010000100110110010100100100111000011000010101101000010010000010001101011100000010011110001100010111001110001100110101011110100111101011000010001001100001111010010011101001000001111001001011001110100110010011011111011001010111110001110001010001010011010011000000101110011000100111101101011100001111011000010111010100101100111101000111000111010111100100010000100101010111101000101010001110111010110111011100011000100011010111101010111101001111010101111000111100000111110100000011111000101100111101001100101011110100010010010011001011110000110100010101011101110110010100100001101100011110101110000011011111110001010111110010001101010100100101010110001101100000011010000110000111010101000101011110100100111110000010100101010110011101000100110100111100000100000110011101111001101011100000000110111010101111010010110001010101110011011010100001101010111010011110110100110010001111001010100101100101110110111110001010110100010011110010011111010010011001111010101011110110111101000000110100111111000011011110111010110100110100001010000001010011000011001100011011100111100000011111011101011011001000100010111011001100001010011011011011111000110000000100001110000101010101010010011101101100000110101000100011000100000101001011011110001110100110111111110000010011101001100110100000100100011011010101110110011110100000010001001100011110011001101011000101001001110000000011100101000000111010101100101010001011001010110000111100100111000000111101010100001010101110000010000110001110000100111101100000111110000001011110101001000111110110111100010011011101010101011111110010100010110101111100010011001110110001001100011110101101000001010111001101111001101101101110101110100011101110000001110111111011110001100000011001100001110111010010111001001101111100010110010000001101011010111100000011111001111011000001111000100100001100110100010010100010111100001110100001100111100000110101110001011000101010111001101111010100010110011011111010010110110110100011000001110110110000000011111101110111000111001011010100111000001000100000100011110000101000101101110100011001111000100011100000011011010101111001001111001100101111110100011011010001111000110001001010001011001101110000011011010101101011101011011011100000101101010111101001001000101101101011010010011101111010011100010100000001011101001011100110010110111101001110001111011010110100001111001000011101100011110111100111111100010100100011001100100101001101010000000010111010000011000010001110111110111101111111010000000001111000100001000010101000100111111111111011011101111101110010001011001011000101110111101100101110011011000011000110101100111101010111001110000000011000011101111001000111110000111111001111010101101000110111010111110011111111001000101111110010110001001111111000001100100000101000110001000001010100010011101011110101000110111100001110101100111010101011001011100101000011111111001011111100110000000001101001111100000001110101000010101001100111010101110000100100101110001111100101100100110100100101000110011000111000010001011011110001111001000010111011111000111010001000101101000110010000010101101101010010101010110110000110010100111010000100001011100011000111101011010010011100001100011010010101000111000001111010101011100000110000111110101110111010100001111110010101111000100001110011011010100001011110100111010010110011010101110001001001100111110010101000011110001001001100001010101101111001011100101110111001110011001111101111010000110011010111000110111100000110100011111011110001010111011010100010101000001101010111001001110010111101010010100100001110011001000011111000011010101101111101000001101110111010111010110111011101111001110011011010000110000111100111011001111010110110010111101010010101000110000101001110010010101101001011101001001010000001001010000001100011111101001011100110000001001010010110101010000111000010011110110110010000110011010010101010111110010010010000101011000110001111000010011001111110100011001101001011000110111110111001100101100000000011101001111110110000010111001101010110100111011000101110110100001001100010101000101000110101101101110000111100101011000010111010010110010010010000111101110000000111011111011101111010001111110010100110111001000111011110000011000000111111010101011111011111000101010010100000010011011101001111111011101101011011101010011111100011000000111111100001011110010100011111110000000010110000010000001111110111001110111001111111101101111101001010111100111100010101110011010100010110010100000111101100110011111111011110010001111000001000011000000010100000000000010101110111010110001100000111011010000001100100110111010001001011000000011110110111101110000001111001010001000101011110000011011111100110001110011100010010011100101110010111110001001011001001110101100100100100000001101000001111011011100011111101010001010010011001111100011011011110111011001000101101110101110100100001010110010110111100110010110000110111010111100110110111110010001011101001000011011010001011111111010100101001010101000001000111000111001000010100001010001100011010101001100111101111010010011011100100010110110011110011110110010101101110101011010111101111110110110010101111101110110100100001011111000010111111011001000000000111011101100000100001010110001110100100111010100101010110011011011010010011101111100111111110111100010101100001111101010101000010011001000101011110101101010011100101001100110111011000011011000110110011001101111111110101011100000000010011111111000101110001100000111000001011110001001100011010110010111001110111101111011111101000001000110111000001001111011111001110010100000111111010011101100010001111010100100111000001000110011010101110001100100001000010111110110100101000011111010010100101100100101101010111110011011011010100110110111011010110010111100111111100001100100110111010111101001101001101101111010101001110100101110001100010011010000000101010111100001010001001010110011001110011111101111010110100111110001110111001100000011001000100111001110110001000001010001100111111011110000101100000010111000001111001111000111010110111011110101011111001001101001000100111110000001000100111110000101000101110000101110010001010110011001111100101101011011011011100111010110011011000100001001100001011001011000011001100110000100011010111101101101101110111011101101011011110010010010010001010111100101000010001011100000111100010111100100100100100011011000010010111110110101110101110110011011011100111101110100110010010011101000000110100110010001100010111011110001000111011001111010101111000011010000101001110100001100110110010011110101010010000011110111100010010010000000111101001001101111001110101111000010101111001010111000101010010011010001111110110110010111000100011000100111011111111101001111101101010110011101101000010010011101100011011110111111010101110110011010001011011100011111011001010110110110101100001001111000100111010010001110100011001111000011111111001100111011010110001001110100010011001001010000111010100001001001110001101000111110111001100000100001010010001010010101001111101001000110100010101011001110110110010110101001100110111110100100001011001001000101001000111000001101001000001101011111010110010011010011100011011001001000111111010011000111101011100010000100101001101111000111100011001100011110110010011110100011101110001101110010010000011101011000010110000010101000000111011101100110101000000111110000000010010110000010101100001101000001100101000000010111001100001011000011001101000000101100010100111001111010001101110011011010101001110010010010000100001110111100110110111111110001111101010111101110100111111111100110101011101101111100111010010110001100011100010010000001010101001001000110111111100111100101110001000001010001101111101000110011111100011010101100000101001000010110001011000010101111001011000010101001101000000111100100110001100110011100111000110101011000001011100100111001101101011111000111110001100110000011100101010101010010010000101001111001101110010110011100000111000010110000001111101010010100010110110001100101101000111101010100000001010011000000010100000001011111000111000111010000110010101010010111001111000010000001111101101111011111101100101111001000101101010111110000100010001111111001111000010010111101110110000001000010101111101111001001111110110110000000101011111000010001110000110010010101000000101100101110011110001111011101101000010111111100010111110001110101011001100001101100101000101010000001010001001111010011100100111100111110010001010101001100111000000110000011101010011000000100001000111110010101001110000011001001000101110001110011011100000010001011101111101001110000101011111100111001000101000101110110010101001011010010001101110011001110100010101001011001001010100000000000100001001100001100110111010100011100110100011111011010111010101001110010000111010100000010010111110000111010000111000111011000001000000000111000111011110001000001000101100010101111010110001101101001100010001110101001011000001110111001111111100011001100101100110001101010100000100011010001001110000111000100100001000000100100011000010001110111010111111100000010000110001101011110100000101000101000011011100001000110000100001110110111001101011011011101100100101101001101100010000111010100001000001011110010010010110110111101100100101000001010110101101110110011011101100010111110111001010001100110100010100110111100000011010110001101110011101100101100011100101011110111000111100111000000010011000010000010111010001100100010110111010111011011000011110011100111001010100111110010110010011011000011011000101110010111011110010100111101100010110110111100101000001101001000101000011110100010110011000100000010101110000001110111111011101110001010111110111000011100001000100111101100101010100110111110111010100011010000000010110001110110101000001111110001101101000110000011101011101000101100111000111011000110111111111100000011100000010111110001000001101100101110000001011010001111111110011110110011111110000001011100110001101000000111101100111000111111011000111000100000100100110001110010001100100100010100000011110010010111001111111101010110011010001000011010111111101001011000110001111110001101100100011001000111100111111011011111011110110111011011001001010010110101000101110100100111000010000100110000000000111000001001111011100010000111010000010000110101100001101010111001110010001010100110101010110011010001010011111110010111010111101110110000100110000100100100000100100001000111010101011001110010101101100001000001101011101110111101111101100001000010110101010000010101001000001011101010001101110111010101101101111000010111100101111011011101000100000010111111111011000101000011110101000011010110010110110000100000001001101100101001011110110110001110000101001101010001100011001110101111001100111101010110110110011000101110100111111010010011100011100110101000011100101110110100111100110100100000101011110011010000111110000111010011010001111101001001010010001111111101111110110000010100010010011111111110111000001011110011101011001110001110101111010001111011010000010101011111010110100001100110110101110101001010000111100101000111010001101100010110100110111111011010101100011000000001101111001101101011101111110110111110010100100111011000101000111011100101111001101101111100000011011001001100100111101110101101111010101000010111110101001101010111001101100101001100100000100000110001010111110011111110001101111001010111110010100010110100001100011101010010011011101010110111101000000110000100011000010111110001001100011001101001111000001110111010111100111111000001101111100100110001110011010111000010000111101110101101111001110011000100010001011110000011101110101101010011011110101001011101100011111001101101000111100001111000001110101001101001100001001010101010001000111110010000010100000100010000101011100010111000101010001110000110000000101000111101101000110101010100010110000111010100001111000111000001111010110110100101001000111000101001111001000100011000111100010010001000010111111101000111101001110110111100111111111111000111101110000110000110100000101100001101110010010100001001010101011101101001111100111111000101000110011001000101111111001101101001010010010110011001011110010011010001001100001010101011110110001010101101001011101000011011011000011001011010001111010100000000111010000110011011100010100110011000001100010010101000000010000101001111001101010110100010101001001011101010011101100001100001000101101011001100010000110010000101111111101100001111101010110111101010000000001100111110000111011101100000101100001111100001110111001111110011011011010100100100101001000000111010111000010100101001000001110100001000100101111110111011110100100000011100111110101011011100101101101101111011001011111001001101010010010111001111010101101001000011111100101101101111000010000110000101100101010011111011100110001001000001111110111010111000110101001010001001111010000001011011110011001101100000111101100011011111100011110010001101010110000011000101001001111111010110000001010101001110001011101111010001100010110100011100010100011010011010011011011000001111001001001001100011100110110000010101011110001010011011010010111010001011110100111000000000001000001001000001101001010101111000111111011110101011010111100101001011011110100011000100101110001101100101111101010101001101001011111011000111110101001010111011101110100101111110010011011011101111101111001100011010010000101011000001111111001010010101010010010101001011100100001000100101110001100010101010110000101111001010101000100111101001100110110101100111001010101110010001111101111101101101000111010100000110000101011111010110001111101110101011011001000011000100001000001010010111000110101100001001011010100101100100011111100010011010011101110001001011010101000011111010010101011010100110110000100101011010010010111100100111111010101011111101001111101010010100110110011101100011100101011010111101010011110111111111100101110110100100001010110001111010010101011001000000101011111110110110100001000000110101111111011111010001111001110100000010000011110011111010100010110111111011001110001000101011100110100011111111110000110011111110010010011111001101001101111100000101010100010011100100010001101111000000100111011001011011001010100101010011001010110000000101100000001011001001111011001111101110010101101101111100100010011110001110110000100101101100001111111101110101000001111111000000100010100001110001100010100111011100101101000011000111101000001101001000000011001110111010011110000101011110101110011001111001000110000110110101010000010100100001110000111000110110010011111100001100011001110101001101011101100010101000010110101000010010000100001011100100011010100010001111111011101011100001000101000101110011000110110110000101011100110000101000111111110010100000101010101001101111000111011100100100110100011101110000010011001001010010111111001010101111010111100010001110110000011110010111011010000001100001110101010101010111111100011111001011000011000100000101111110000000101001111001011101010001000110001101111011110010110010110010101011111100010010010111110110001001111111011011101011001001101101011101101001110010100001010011100001111101010111110000111001011110110001110001000011101101101101001010001010111101010010111000100010100001110101110101101000001001001101001101101010110010111111000010001010011111110010010110101100011101101001110001111111100011001101111101000111101110000100101101110111110001011010010011110011000101011000110011111111010000001011010110101011001010001111000011001110101101011101010100000100101101101001111010011010111100001000100110010001010100010011010110110001100100011011011111001110111100011000010001000100101110001110101101111100111101011001000011010110000011101101111111001000010001101011101110001001001011000001001001011000011000100011010110110001101100011010010100100001101110111101110101011010010101111011011110101111011100001011100010110010011111100010000100111011011111011101010010100000111110110010111111110010011011111010001001111001111101000110100000001011010011010001001111100110000001001010011111111011111111011100000110111110000000100110100100011111111100101111110101000011110011101110101101001111100011001001100000010101101010101100101000010110010011010011101110101011000111100001110001000111111000000101111110100011101111111011011111011110011110010011000011101110011000110111111110111110001110001001110101110010011111000010010101011101111000110111010001100110100011110110000010001001001000100000001011001101000011010101010001000011001011100101101110110000011001001111000000001001101011001100010001101000000111011110110101111001011101111001110100011101100010110110111001110100000111111001101000011011001000000111110100100010010110011000011000011010000111101011100010001000011000101000010001010101111100011100110001010111101110010101011011001001101000111011111011110011010101101000010000110001100001101110001100011101011010010101010110101011010011100011000001001111111111000101011101011101100100001001011111100111011100100001000010001001111001010110010001100000111111111000011101011001101100110111111101111000111010000011100101101010001011000011100010111111100100101011101111110100100100000010110100101011010111110000111001110111101111110100111111110000010110100000001101000100100000011011011000110111101100011101010100011110011101100011011001111000000000110000011100100011000011011011111000010111110101111011011001011100100010110101011111100110001101110110010110010101001010000010111001100100000010101100110111111101110011111100100110100110000111110100000001011110001000100100010011100001101001100010001000000011001101010001000011100001000100111010011111010111011011000111001111100011110010100111011101000000100100111111111101010001100001001011101011011010111111011011011011010111001111011110100001010010101010011000011100010101111101101111100010000100100001110000110100010010011111100111111110100111001001011011100010101110000010001000001010000100111011011011011101100011000100011001100100111000110010000001101011101011101011001111001100110110100110010001001010000010001100001111111010000000100010011001010111110110011101111110100001011110101011101101001110110010111001100101101100111101101100000010100011011110001110110101101000110110111010010010001011011100111100010001010000111100010110110110110010100100110000110010011010100101101001001001100100111111100001000100000010101010101110110101100001110001010001011001101101110100011111000000010010110001001110010010110111111100011100111011001101101111000000000111100110100001010101011111100011011101010001110010001010101101011010011000100000011101001000110011000010011101110000111011011100010100000110001100111001100101111111011001001000010101111111010111000101111001010000111010011111110000101000000100101010110011100011110001001001100011001101101100010011100110001111110100011010101011011001100010100101001000011011011011011000110001001010010001110111011011101100101100010111100011101110011111001101011010011111110101001000011001010011100000011001010000011011011001000000111110011011001001001111000111111110111101010101111101010000110000010100011111001010000101101011110011110101001101100011001100011101111001110010101001110000000000101000010000111011011110010110010010010111100111111000011110011110000011100010101011010001100001101100000110101011001010011000010011001011100001001110001011110001010000001111000011001110001010111000111111001011011011000100010011000110110010100111010010101101011010110000010001011001100100001010000111000111010000111000111001010010001100111000110000000000100111001111000101000101011001010010101110010110001100000101110101110001000110000011100011111100001011110111100100000111101100010101010101110011100100101111101100011100110101100001011111000000111111111001100001000000101100110101111111000110110110001001111110010000111111001000101100011010110100111001100010010010110011111111101011110110000100000001110110111010100011011001011111110000100100101111111000101000100011101111010001011111011110111001010010000100011001101001100100111110010111000000111110001000011000011111001011000100111101010100110101001000111010010111101100010011011001000000010111111110100101100110101001001101001010110111111001101000000001111100110111111011101111000111100000000000111101011101100101111101001100111100101110000111010110000111100011010010101111011000101011010011100010111101000010101000101001001111010111010111110100000101010011110110100010100011010100110100010011101000100000101001111001111100111110000101011000100011110001011101010101101100101111001100100101111101011111011111110010011000100100010110001011000101101010111011101000001110011110011110000011110010011100100011001011111000011111110111001000011000101000001110100010100101101100111011000110110011101110111000100110100100101010110011111110001111101001010000001101001110110101111100011000000101110000110111111101001001111011100101110001000100100101100001001101101010000110000100111110010110000011001110010010101001001000001111111100011011010011101110110110010000001001011001000011100001011110000111011011101111010001011010010001000100000110111110010001111111000010000110100111010010101101101010110001000111101010010111001111010011111100101100111111101011000101010111001010101100101010100000111100101101101001100110010110000010010011000110100101100010110001101010010001001101101000110001110101010001011010100100101000011010011100111101110111101110100001101101110100111011101010110111001101001011110100000101011110001000111000110001011111000011110001111000110101000001111000101010111101101100101111101000100001010111011110001101000011110111101010001000100111110111010000000101100100100001010100111001101000000010111010110101011100001010100111101100111000111101111101110111100001100101110000011100011011001011101001101101111000001111000111000011001001001001100100001000111010110100010111000101001110110110111000100110100010110111001011110010101101000110110101010100101011010110000011111001011001110001100111110000100110111000100110101111011001110101111011100101110000000100100000010001100111101101100100111001110101011000100100110011110001110101101100001000010101011110100010101000001100110110000000100111000001001000001010100101010010110100010100101000111101010110110110101101001000111000111101100001011000100001000000111101000100010111010100100101101111101110101111110000100111111111101111100110111001001100101100100000100000101111011110100111110100111000111100000111111110100100101110000110101010000010100101100001110100110101001000101101000000011110110000001011010100111011110010010001101010100100000011111011010000010110000101010011011111101110110000110100111010110111100000101110100010101100110100001111001111110110000100001100010100001100111010011001000111000111011101010010011111101110000010111000100001110010001001011000000011110111100000101100110010000111110111000001101111111001000111011111001101111011010010000000100010011100100000001001000001111110001100110001010101000011011010011111101101111110101001110000111001100000111111010110111000100000101010001001110001100000100011011010101000101001100000110001101111110011110001111110110111101110101001001100001000001101100010100110001100011101000011111010001001111000111101100100001100111111001101011111000010101111011010001101001110001111010101010011111101111001110001000001000001000100111011011111001001001101110110011011011110111100001000010101100111010011011000101111000110011100000100101110000000110100110000010010010100001101010110001110111011000011010001010110111000011101001100011101110000001000010001011111110000101010000010001001101000000101011001100111111101100000010000010100101111001100010100001010010000010100010010101111001101001011110101001000010100001001111001010010000100110001100100010000111011010010111100100101001110010111011111001101110100011101101111000111111011011011011001001110000001110111111001101001100000000000101100001000100001010000101001110000110011111101011010111000011100111111000000110111110010111010001001010001001000001000001000111000001001000101101000110010011110111100010011001011110100111100101010010110011000110101010011011110000000011000001011001000101011001110111100010010110110111110010110001111111101011000000011101000011101111111011100101100101011000101100111110111010101111111101010100010010011000000000000100101100100110110011010101100011100100000110101011001100000001101010101101100100010000111010010100110100101111000000000001110111111110101011100011000110000111011111100111101000100011011110111010111100110000100011111110010010110110010101011110011101010011000011011001001011101001010101000100100111110001010011001000100001001101111110010010011001101101011001101101000011011010000011111001010001111111001011110000111000011100110100110100111011111001001110110001101011000001111100000110110010011110100100001000100111100100111110010100111100001110100011111110111011100001011001101010001110101000100000001000111001001101110101111000111101111010100010011110011101101001010000110010001000101111111000010111101111010100001110010111010100110001001100101100111001011111100101000010000000101011000001100110100000001110110100110100000111000001100100011110111011110010011100000101001010111101101010011110100000011100110111111111100110000001011100011111111001100011001011011101001001100110101001101111110110000101101110111010001111010001010101101001110000110010101111111101110110000100101011011101000101011111001101000001010111110111000100101001110100010101110100101000001010001000000100110011011010110111011110011101001011101010000111100010100111001111101001100101111111000111001000101110000110000111100001101010011001110000111000010010001100010001010000011011101101100111110011000110101111100110101100101000101000001011011101101111111000011110101010001110111000101010111111011101110001000011101011101001110110100010100110110111111011010000100010111010110011110000111010001011001100101100101001100010010111111101010100100000001010111100001011001001111010000110010100001101100011110011010101110001000110101110110010110000000010101000100010011101101001010001001011010011001101011100111100011000111000101111111010011010110001100010111110110010110111000100100001001110100101111100011001011010101110011100111010101011010100011101010000010010111001100011100011101110110111000010011111010011000111010101001110110111100010011100011011101111011110000110100011011110011000010001011101011101010111011011101010001011111111100011010111001000000001010100111010000001111011101000100001100110110000010111110101010000000111100011111111001001100101001010111000011111010011110000101010000100000101100110000111111000010101000001011010101111000000110001001110110001001111100011000111010100000101110100100111011000101010001101101001010100011111001101001001000011010011111101100011110010011111110011101010000111101010001001101101100001110010111011011110101100110000111000100100110100101110110101101100101111101011110101100100000011100000010111111111100111001010100100001111010001111101110000100111101000111000100000010101001100110011001111101110011110101011011001010110001001010100011111100111010010110000001101011000111011010100010011110111000000100000010101011010101101010000011001111101001110110011100111010110100100110010001111010110011111101000011111100000001010110111001110110100110001111000111101101001010111000111000101110111101101111000110011101010110111010010010001010101100111100101001001111100010000001101010010101010111110001011000010110100101100001001000010001111001001101001100010011100010000000010001111010110001010001010111101101111110000111011100010111010100100110011111100011000100100000011101010001110011111001100111111011110010001011000100011101111010100100111110111000011010001110000110011111100001001100101101101111010110010100100110100010101101111011000111101101011100001010000111001100101001111110110011010111101101101011011110010000010101110011010001000010111010011001010001110010111000100111110010010001111010110000110111110101010011010110011011011100100100111100111001101111010101001110111011111010101100110111111011100001111100110011001000011101101101010001001110011111110110001011011110010110111001011100110011010001010110110000111000100100011110011111000110111011110101100011100100100100011001101000010000110101000011000100100111000011100110111010011011011010001010101110011010010011001110111101100111110001111010010000111110110101011110101111001011101000001010100101111100101110000010110110111010111001100101000111111011110000110001100101000010110111010011011001001100011011111101101110111011001010001100111110110001110110000101001010000001111110100101001111100111111100101111101011000101011101100001110001101110011110111010101001110110101101101111011000001110010010010100111110101110011010100000011000010011010011010111111001001100111110011101011110100100110111101100000010001000110010100001110110011100000101010101110011110001110101100010011101101100011011010000000110010001011010011111111000010101101110001110010110000110111111010011000111010111001011100101110111100100110101100000000111010110011010100010000001100011111111100100101011100000110111101101100101000101111100000111010101011111110010001101000010100100010000000101010111111011001100100000100100111001100000101101100001000101100111001101111100111001100010001101010101011001010101110110010010100001100111100011100111000010100111001010101011000000101111111010111110011100001110011010001010110000111110110100001010101011101011101100111101010010010101110011001011010110000101001011010110001100101100110100101000110100010100011010001111100110000110101101101111100011000010100001101011110110001100010011000111011011010011100101010100100001100111000010100010100000011001110110010101111000000000010000000000111000001000110111100110000010000001111011101001101001110011110100110010011101101101111111001011011011100101101101011100001001010001001001100100011100001110111111001000111000000110010101010101100000000000010101111100010000010000100111111000101101001011011000110100010110110100111001100011011101100100001010100001001100111101011001011000111110101111100011000010001101010101000000001001010110101101001111100110001011101001000001000000010100001010001111000100000000110010100000010101010100010100010001000010101010010110101010011010100011100001001110001101001100001000111000000001101110110100110101010100101010100110001100011001110001111000000010100111000000101010000111100100100101100101000011101111000110100101111011101010110010000111001110101001101001100000110010100000001111010001101011011011010100111011100001000011011001101010101010101100011100000100001101110111100111010100100000000100011111011111000000100100001111011000010111011100111100011011101111101110011000111111111111101010110000010001000001000110110111101011001000100011110101001001001001010110100110001010101111101101100101000001101110011001101011001001111111001010110111110011011010111100100100010000100110110001101001000110010010010011000111000001011011011000111000110110111011111001010111000010011000000011000111101100111100001111010110101110010111110110011000011110011010010001101101000110111010111010111100001101001000000101001100111001011101011111001000110110001110010111010010001111110100001111011100101011110010001010100101101110110101010000101100111101011100111100111001000011111111010011011000000001101010000110111111000010011011111111111110101111000110111001001100111001101110100010110111100111011010001101110100111011111001111111010001001011110101011100101110011101001010010010001001010100111110110101011101001001110110011010110011010000000111100111100100111101100110000011100010111010100101010001101001100111010111110111010001011100010100011010010010010110111101110010001010011111110100111000111011100111011000001000010011010010011111101110111110100111011110011010111001110110100110110011111010110111101011111111010011010100111110111101111010010001000100100111111001100001110100000111001001011111000110110011001010100110101010001111101010000000101111101001100110000111010001000101111111111001011001001000010101010001001001001111111111001111001101011100001111001010111110010100111010110110110011000101000111011100100011100101001011010011101110101000110001101111001110010011110110110110110010101100111101010111110110001010010100001101011111100000001000010111000000010110111000001100110111111011010000100100100001010001010010110110101001111101101100101110110011100100000010000101011101110001010000011001010101001000101101010110111000100100111000011011000101110011011111010001000110100100010011110100000000111111110101010000111010101101011110010001110101101111110111101110011101010111110111001010100010010001000110010011111110101100100001000010001111001001000010110000110011001001010010101101111000011010011011110111000011001000001011110100010110010100101101011111010000001111101111111001111110101101000011001110000111011011100110100100110110110010010011110010010101001111010001100011000100000000000001000101000101110010110101001101111000001000011010000100111100111010111111100111111101000111100001101101011010111010101011011000110011000111100110110101000111001110000011101000100011011000101111111001101100101101111111101011100010100011010001111100011000010010010010101100001010001001110111110110010000001100100110111011011111110011011001001011011110101000000001011110100111000011100001001010010001011111101011100100000001111010111101111111010100111001100000011011101101011110001001010101000011111011101100000010100100101111100010011110110101110010010011111100111010110101011111011000010011111001010000111101001101111111110011100100010100000001111000001010110000011011010010011010100110100110011001100111111001000000001011001101111000011000000000011101010110011100011110111001111111000011010011000011101011001000100011011111010100101100101100101111110110011100000001001011101001000101010010101110011000000111101110010011010110001110000001111011101100010000110110101000001010011000000100101010010100000000100110011001010100010110111101101100101100010011101001111100000010011101010110110101101111111111100010110101110000010011101110101111010011010111111110111101110110001010011110100011010011010100111010111011111110100111011011110000111111010101100101101011000100001111110001011110000100100110111000100101110111010011111110001101100101001111111100110110001010110110001101000100111111100110000000100111111001010010111001011101001001001010000010010100100110011100000011001010000010011100010000010001100011010101000000100111000111101001011010010111000101111101011100011110101101100011110100011000100001001011110011000101100010111110101100000100011001110110000100101010100000101111100011101110001010101001000101010100000101000001010010100011001001011101101001000100010010000101100010101010101001101010010000110010011111110110001100000110101110111000001110100000111100010010101100110110010001110111100111101100001010000111001011010101000111001010000001101100111001110110010101110011000110000001000111101101000100010101101001111011000011110010000101101001011100011111100110100001110001000110100100011010110011010100100010010000000111000001110000111101111100110000000001000111100010001100111100000010010110011000111100101110000010111011011011001100010010010111010101110000100110111001000001111010111101110011100101011111000111110010010001000110110110011100000111000111110000111101101100001101110011111011110110001100111000000100101010111110101000010101001100010111010100010100001011010010101001001000010000110100010111110011110010010111001101101100011101000011111101101100011000110111001111101011111010110010011110100010110001011001011110110110110000010000010101000100011111100110110001101100010011111001001110010011000100001110101100100111011000110000010011101000100010010110111001011100110100000110111111111000111101101111000110010100001111110111000011000011111010100010001011010101101011101011111100100010100100001111011001010000001010101010100000111011010011101010001111100001000111110000111000101011010000100000110100110111000110010100000011011101100001101100101101011001100111011011111010100110100000011111101001001101110010001011010010011001101000100000101111110100101100001111000011100000110011110101010110000100010011110001000010000101101101010100010100110001110100000101001101111001000110110010010000100000111111101110100100111011101010111000000001111011000100000111001010111101010001011001101101110000010011001111010111001111011010000001110010100001010001011110001111110100011100001000111001010101001111010101110100010110100111111011000111101110000000011111010100100100110000010101010110011111001010011001011001111111010001011101101110000101001111100110110010111110110101000000101000110111110111100101001100101110010011111111001111001101101001110000100000000100011110110100001100010100000101010101011101101011110101001101011000111011000101100000011010011011111100101000011111100001100010100110101110110011000111101111100010111010110001001111101000111110010001011011100100110111000001000000110001001101001101011010000001100001011011110101101110001010001001010100101010110110110010001001010010001000100100101100100100110011010011111110111011111100100110101011100001100000001101111001111010011111110001000001111000101111010110000011001011000111101001111001110000101100010011010010100010001101110010111000010010101010100010111100101001101110110101010011011101000100111010101100110111000010100001110010000010110010111010001111111010111010100110001010001000100110010000110100100110100011001000100001000100000000100111100110100100100110001110101010000001000000110101010111011110101000101111101101101001111001101001111001111001100011011101100010001110011001001100100100011011111001000001110010011101000101001011001101111010001111001011010111011101110000000101111111010011100101111101010011010001101111100011110100111111100111111011001011110011101110000110000000100110101101001000000010011100001111101110110110001111010001011110000001101111010110010001001111110010110100101110111101001001100000010101101011111011100001000110101111111100100001011110010010011110010100100110001100011110100101101101011111111011111010111101111000001010101110001111011100010001100111011111100010001101100010110101001101111010010111101110010110100110011100101100111110100010111011010100000001101111010011101111110000000110111001100110111111010111100111000111001001011001100000011000000010110110011111101011010001100111001101010000101101110000011000110111011100100011111011100000110010011011001011101010100000111001001101101001010011000101011101111010010000101001001001111110111001000100011010111010110100111111000101010100011111111111010010110010100010100101010000110011000001010000010111101010111100110010001001000111010111001010001111111100110111010001001100111001001110110001111100010101111101111101111101100110000010001110011011111111100101000010110001010011110110011000000101101101101100110110010110011111010100011010101011000100100011100110110000010101000111110000001111111101001011110010011001001100011000100011001100100011100011111111100000110011100001000100100010100100100011111100011100100001100001011110110010010111111110110000110001110010101000011000111110110101001001000101100110001011000110001111110010110000011011000100110010101011101011111000001111100100110011101101000011110101111011000010000010110101101100111010101010111011100010111100011010001001100000101010001001011000011000000110010011100011000010010111110100010110110011100011001111001101111011011000101001010111000100111101100110001000100001101010000111011111001010001101010010101101110010010110110101110101110010101100100100001111011111001111111001111110111001100101001011010110111101111011100010100111100010001100100000001000010010011111101011111010111000101001011101010111011010111101100011011110011001011111111111111011010101101100001110100101110011111011100111111110010110010100110010100001101100011010011010001101010001101111100101111010100000110111100111110010001010110000100100100110100010100100110010000011111010011001001110111011110100101111101111111001101011110100101110000101010101100101011010010111010010010011110001000101000111000110000101000001111110111010001110010011001000101000110001010110001110001010000111001000110011110101111001110000011111110111000110000001100011100010111101000101100111011001010111001100100010011010100111111110011101011111010000010010010010001000100111000100110111111011101011110100001000101001100011100111011100010001010101000000011001111011010011100100111000110010110101110111000110100001111101111001000101101100100001010110100001001101001010000010001101010001001001000110111011000010101111110011010110010111110110010100100111000001011100110110111010111001010101111001011110000001010101110100010100110010001101110000010111111110001000001110010000111001101010010111110010110111001101001001111100000111101000011011111110010101101010101000010001100110100001101100101000100010100101111011001011001110101111001110111010111001011111101001111001110001111011001001011010111111010100000100111101001100010010110101110110101001111001111100101010100111011011100001011100100101110100100010111010111001111001110010111001000111001010001000011011100000110101011001000001000111100111010011111001000100111111100100111111110101101100101111001110011010100010111010101100011101111111110000001011000001110001011110111000101110100001001001100111100011111001110010100111000000111011010111011001001011101101100011000010000100100111011111011110001100000110110010011101001011100111011110101111101011000110000000001111011101101010111011111101100110111010100010000100101001000100111110111101100101011101001110111010000101001011001111011001100101100000000011110111011100111100000100001110101011010111101100110100000000010010111101111111010101010110010111001011100111001100110001011101101110000010001111011111111111110000111000011101000100011010001100010101000000111111001111100111100110101101001001000110000000101000101100000111001100110110011010001100110011111000010101011000101010010010110001010011110111111101100010101000001010100001110110101011001001110111001001100000000110001011100100010110110000101011100110001000101010100000100010110110111101100011001111101010110011101100111000011001111101011101110100110101010010111101000001000010101111101000011100011011110010010110101101010100101110101100001011000100000001001001111000100101010010001000001111100100110111000001011100100010110110111011000111110001011111011110100010101101001000110101100011101110000110101110111110000011010011001110111101011110000001011001100001010001011111101111101100111001011111100100011001001011000010010111111111001011100110101001011000101100111101101101100011101010011100010010101010001001011110000100110110000010001010111000101111101110011000001010101011110111000010001110000100011111001011101000000110110001011101001011110110110000010001010000001011111101110010010000111011110110111001111100101000000000100110111010100011100101001011100001101000101100100101010101101100110111101000101110001000111010100111100000010011110110001011100000110010100110010001001111110110000001111001000010011011010110111010000101010111011010111100110101101111110111001001010110001011001000000000110000010011011101001110001000011111011111000101101100100100100100110100010110101011010100111000101101101111110000011100001111010100100001100001100100000101110011110011100111010011000110010011111010000111100111100111111111100011010010000010110011111100110110111100101100011111010101101110101111111011000010001011001010110001111111011111111011111101110111111010110101100000000000110010000000011111100010001110011101001100000000001101011100101101110001010010101101011110011000111011011111000101100001010001110101110111000001001100101000011111101110111101011110110110010000010010010110010001110010001010011010101011001011100100101110100001011101101110000000010111001110011000011110110101110011011001111111001111010111100111000000000001100110001001000001011011100000000010101110010011011110000101100000011101101101010001110111101111111101011101001110011001111001111001011100010110000010010011100001011000001100001111000100011101101110101100011101111110111000001001111110110011111010010011010011110101000010000111110111001010011100011100100111111010001101110001110101000010011001101011000111100010000001110110000111011111100001101010000100001111000010010000000110010011000000111001110011110100001111001111010010001010000110010111000101011010000010001001110110000100000111100101101101001011001101110001110010100101000111010111000010111100111111101110110011000010111010111111110010100111111011101100111100010001100101011111010110011100101000010111000101101011011011111001101010110111010110111010000111100010011000110101100101011010001001111011111010100110100110011011010010000100010101010000100101001011011110010010100010010001010110001111101110100100011111110010111010010011111000111111111111111010111101111111011111001010010011111110111001001110100011001110000100010101000011001111111010011000101010010010100011101011100100111101010101101000110000111111000101010000101110111000010011101000111010111101101110010001011101111100011001111001000001000001101010010010101000101101111100110000110011001110110011000110110100100111011111110111010010000001001011110101101100110111011101110101111100010110110110101000001010010110101101011000011110000011010111100110111011001010011111110010011110011101001110100000110010001111101110110010001000011100010000001011000111011010111000000010011110101001100010110101110111111000110011011110101011001111000010110110001101000001100100110111000101000001011101001001111011110110000111010111110010001001011011010100010111001100100100010001100110000100110110001001011101001111110101010010011111101110000001100110001001010100111000110111111011110111110000101110001001010110011100000101111011000100111101000001100001111111100001101100001100001110001100110101101011101010101001011010111101111110011110001101001110100111011111110110110111000110001110011010110001101001101111100000011001101001110100010010101101100101010110101001100011101100101000000010010011010111010011111100010101101101001011111111100000011101001100100110001010001011111100101110101110110010011000011110111101111100111011011001101001010010011101111101010111111110000111100100111010010000100110111010011011111101010101101010000001000110000000001000010011110010100100100101010110101001000001101000100101001010001010000110011111101101110111100110011101100011100110000011011001010000000001000100001001000001000110101010110011010110101100111001101110101111101100011110001010111100111110111110010001100111001010111001000001011001110110001011110011011000001111111010010101010100010011011111000100010110010111010111010100011000001010010100100010011100100001100000010011010100001001010010010010010000010110100000011010001001100010100011101111110000001000011111101000101101100011000000011110101100110010000111110010001011101100010001100011000010001001100001000101111010111000000110011010100011101110010101100110011011010100110100110010000100000100101000100101110101100010111011111000101100011101110001000110110000100000100011101000110011010001010011010010010101001001011110100101000001110000111100010001110111100011000111001101010001111011100111100011001011110100000010011101011101011101011011001111010110100001000110110101111100011100010100111000000110100101111101000111111000011001011000011111010010001111101001011011111110001110011110010000001010000010101110100100000000001011100000100100100010011101010001100001101100001111101010101000001110000110011101101000111110100110001001110000111000001110010010011001000110011000011011100000010100011011000010010001100110001000101100000000001000011110000111100111110011110000110001011110010001011010111110100001110110011011001000010010010011011110111100100110100111001000111010010001110101000001111000001110011011111111100110101010100110111011011000001001111010001000111111001011111100110010101111011010000010111100100111101111010010100100010010110011100100000101111111010100110001110000100111111000001100111101001111100111010001111011101001101011011010011110100101110111111010110010011000001110011010000101110111001000001110101001110100011100111001101001011001110100110101110011001010000110100110011111011000001111000101001111110011001111010000100110101110100011110110101010001001111110001101100110110101010100001100111100100100000011000100110101000110101100101010101101111110001000111101001000001011111110101000111000100110000111100010000101111001000110110010100011000100111111101010110011010000111001001001100111000011110100000000111110000011001100011110010101101100001111001000110110101000100111101111110000011010001100010101110011001011011111101101010001000100101101010001011100101100101001100101010000010011000010011000110110010101110110100111001111000010010010001001110011000000101101001001100111110101111011100001111000110100101011010110111101100111011100010100011000101000010010100111110111010000011100011111110000101010101100101011100101111010101101000011101101001011110111101011100010111111110100110010010101100011111100110100101110011000101000011000111100001010100010000111011000101111101111111011101011100010001111100111111011100100010010000101100011100010011110111100101011101010110100100110011100100100011111101000001010100000111100000100110010010001100110100010001000101111010000101001111100001011101001111010110011011000101111011110110000001011010100100010100110001111111000101010111111101101000001111111001010110111110110010011111010101011111111110010110010001011111110010111101011010111110010101001011010011100100010001111111110011000010001001100010011101011101010011011110001001010011000000110110001101101000010110000011001000111001110100111011111011001111001100100001101111011011011101111001111110001110110100000101000101101111111110110010010001011001110100111001000100000011110000000011111011011001101010001001110000001101100100001100010000010111001101001101000011011000011101000011110110010010010101100100000101101100001110001001000010000101101011001111100110011001000010000010100001000000110000001111101100111101111011001011000010000101010100100010001100010011011110101110011001111111111101010010100100100111110111110100011110010100010111010001001110000000101100110100111101001100100110100000110110111001111000101110011101000010010101010111000010111011101100111010011101101011010001001001101110100100101011101101101001101111101001001100010001111011101111101000000010111100111111101011111100101100000000011110001101011110011100001101010111000010110101011110101010001000001010001111100110011111011010101111111101001100000111011111001110101010110010110010010100011101010010011001011000001101100010001001001000111110000110010101101001000110101010101111001100111000011101011111011001010001011001001010000111110011011101001110010100000110101011100010011110010011101100000000010101001101000111010111111011010101101110100101111110010011101101101110100101101110100101111011011010000100010000000110101101010011111011011001001001111111111101100011110111111010101111001111001100100100100101001001100000100100111111111011101111100111111100011000001101001111111101110111110111011001111101000100001011000011001000100111001100111100000110111100001000001001111101000111100011001011100010000101100101010001010010100010111110010011100101011000111101101011001110100001110001111010111010010010000100100010100000100011111101100101111110001100011110101000111100000001011001100110100110000001000110000110011000000111110010001010000101110011100110101010001000110000100101100010010011101001001010110010001100010111011011101100011101010111011100001000011111001000010000110001100000111011111001000010000011010001100110010001100111111100010000001011011011000011101010111001101101011011100101100100010001010001111100110001010000001110011111010010100100110000100000001011011101100110010111010110010011010010000000100110010011101110010001000101101001100011000111001011011110011111111111000000001100100110010110101011010011001001111101000100100001101100011101010001100011001110101001101100000011111001001110001110001011111001110000010011000011110101011111100010100111101101011011101011100000010110111010010101100101010101010011110111111100111101000110010110000011000101001011001100010011101100011101111000000101100101110011100100001101100111001110110111011000011110010000100000000100010001101111011111010000101111011111011111010001000101101111111110001000011110001110111010001101111001001101001011001001011100111011100000010010100001101111011101111111010100000100001110101101100001111111100110100011101010110010010111111111000110000011011011110011001011001010011111101101001100111100101001110011011001110111011001000000011010001100101011101110101011100011000001100010111000101100000001111011100000011011001001100011101011010101110010001010111110011111101010100011100110110000100000111000100111011110110101111110011001000000101010011101100111110111001011110001101001111111010100001011110101111101100111001001111000001101010000001000110100010000000100101101100000111101001101101100011111000100100000010000010110111111101011011010010010111101111010100100101100110001100100101101011101001010011101101101101000011011111111111100011001010101011111111111001001100100100001111101000110110011011101010011000111000001000101110111011000011011111111101010000111100001010100100110011101111011000100010000001100101001111111100000000000111110110001111010010011111010110001110011100110001000010000001010110010000010111010110010000111000111111011001111101111100000001101111001011011000100100000110101111000110011011111100011001111111001000110100010010100101010101101100110011111100000101011001011101110100110110010000011010101101110110000011111100101000011100001101101111000000000010011001100110011100011100110100000000000110010110010100011011110010011110010110101111011100110001100000001111111011001101001110000110001011011010110011001101001110100100001010101101100100010111001011110101101111001111011101110111010111100110100101110011100011001000111111111010011011001101101101110101100011011010101011101110000011110100111111000110010000001111111111101100010011110111100111110000000000111010010000011011110011111010010101000101000010000001000110100100110010101010010011111110000011000001011000110110000110111100100010010011101111011000111000110001111101011101100110010010101100000101101010110001110000010100100010100101100111011011010100100101111011101000010100111110110001101011010111000110101111000110000010110111110110101001110111100101010111111101011111100111000110001001000000110111010011001000011000110111100111111101001011010111111111000011100000000111001000100011111000001110111011001001110110111010100100001111010000001011111111011011010000010110111110111110100111011000101010101001110111010000100000001101010001110100100111011010000110011110000011101001001011111111000011110000010111001101111100011101101001010011110101000010001101011100010110111100000000101110000110000110000101110000110000111101110101010001010101010011001100111101001100110011111011110011111001001110110011100100010110111001111100011111100100110110000001000111110001101010010110110101000101010111000111100010101010001000100101110100100101110010001001111010001110101000000010001111011100110000001010010101001011001111110110111000101110101100010110000110101100101010011011001111111101000001000100011010111100000110010110110000101111001110010111001011011010001100000010000000101101111111000000010000100001100111100110110001010101010110111101011110111001110010100101000000110111011001010000100100000001111010110010100101010101000110111110111011110100011011101000111101101110010001110011000111101111000110111101111100000111011001111011100010001101100011111110011000100000100100100101100111010010101111111101101000010111011100111000100111110111010100001000101101110001011001110111100110110111010010011110010100000100110110111110000011111010111100110000000110000011010001110010001000100111001111000110111110111101010001101111100110110011010000000001101100001001110011110001011000111100101010111101101001000000010111101010110111100110000010101010001011011111110111111010010100111000000110001000001110101001001100010100011111111111010001011011101001010000100111010100010011111111001010000111100100001111110010000000110011010001101100011110010000110001111000110000101111010101010011010001000111000000100010101001101101101011111110011111101101001101000110011001100101001001100100010010110101110101001100111001000001100000101111011110011111011000001010101100110001110011101011001101101011100001100111100110001110100110000001010101000001000111001110010000100001001010011010000101101011110101000111101100100011000011101000111101110100101011101100011101100110110011010101010110000001011100111100000010000100011000100011110000110010110000010001101111010011100101000110001000110110010001100001111111110010111100010000001011000000011101110010100100111011100101110101000011000100000011111100000010000101110101000011010001011111000111011110110111101111010101000001110000100111100000000101111011111111100110101101111010011111001110101111111000101100010011110001110101110111011011000010001001111001010110111010111101000100111111111101100101110110101001101101010011010110111000000101010111101011000011110111011011001010110011010111100100010111101111010111011000101101101000000000010110010000010110100100100000000110101000100100011110101001111011010001101110100110011000000101100011111000110111110101110101000011100111100001110001010101010111000010001101010100101011100001010001000100000010001101101011101001011001111000011111000000101111110100001111111101001111101000100111110000100001110010111111000101110011000101000110001011111000110000110100001110100001011010111101001110011100010101110110011110110110001000010101011000100111110110010001000101000100000110010011101111010100100011010010010111001110100010010000111111111010110000010110100011111100001100010110100000001110011110001011010111101000010101011111100111011101001111110101001110110101011001000001111100011011101100000011011100010101110001110100001100010011101100101100111111000101100000100001011011010101100001000110010110101110101111010000111011000111101001010110000000111111001111100111110101101011010110111010000011110111110011111101101010011110011111100110001011100000000000111010001000111101011001110111110001011011111001011111011010010110011001111110101010101000010010111110110110000110010111110111111101100011101010111010001000001100101001101000110010001111001010110010110110100011010111001000110100111101111010001100100101001000111100100101011011001100010001011110010101111011011011110010001100101101101001110101111011000101000101110010110001010100111010011010000100111010100001000011001000100100011110111101111000110111011101101001101111011011010100011101111011001011111111101101001011010101111010000111101010101010111101000010110010100101010010000000100101110110010110111100001100010111111001111110010001001111110011101000000100101111010001100011000011101100110010111110011101100110010000000001011000111011010111101101011110011000011111000001110100111110000111101110001110000101111010111110010100010111001011101101001010010101011010011110011001100001011011011111000110100111011110101111100110100011110000011010101010100000010110101100101000110010011101111011011010101101001001011101010111001000111101001000110100100111011010011100000100110011001001001011100010100111110000010001011111011011101111111010111011111110101001000010001010011011010000101101000011110111001111011101101101100100011100100111010111010101110011000010110110011110100111010001111100011000101110111111101101000100110100000110110110000101101010101001100011010011010111110100010111000000001010111000110100001011000010101101001100110101101001110011110100000011100010000111010101101111010110111001010011000111000100011001010001101101001110100111110010000000001000010101000001001011001111111101011100110111111101000100111001110110010000001111001010111100110011011010101110111110010100100101100011111011001001110011101111011000110000110001011001011010011000010111111100000001000110101010000000100110111101010011001001101110100010101110110111101111101011101001101111100011011011101100100100011001000100100101000111110111110100101111101110001010101000110011011010001111011101111000101001100010011100111010101111011010110001110100000001001000100111010110110010111010011110100001110001011101101010101001111110101111111101101010000101010100011000001011010011111100010101001111110100011000101111010101000100100110111011100011110001100111000001000101010100001110011010001000100001111010100101110101111010111010101100000010111111011001110000110111001111001001001111110011001111101111010001100000010101101111011010101010100101001101110100011100110011111100010101011110010010001110101101111101000110010100111001010001100010010011000011110111001110001000010100000110011001000000101010111011010001010101000001111101100101010111011101001111111010101101010001101110111100000011111011111111011010111110111100010110011001101101001000010101000100101111001010000100101001111010111001101111011011010100000000010101000010111100010110101100011010011011111011110001101001000000001100111011101101101000101110010000011101110100100100001100101011110110110100011100100010000101011111110001110000110111011000011110010111010110010011100000000000010011101000110110101110001101111110001110001101010110011100100100000110001101101011010010010000100101110111000100010010010000110101110011010000100111011000010000011011101011001110101000111011110111010011111110100101100011000100111000111001011011010011000011011000000001101110000010011000101111111000100101100001011001100101110100011110100011010000111101101111111110010110101100100111100010110010110001111101111001000001011011001100000101011001010100001111101001111001000000011011011010000100001110101001111010111000111111100011100101111110110101101111111010001111001101101111000011000101010011101100100111111111111000011100010011001001111111011000101110110010010111001011011101101110110101101101100011111010010001101011100110110101001111101111100100111001110001110110000100110111101011101100101101000101010001111100001101110111011011101001010011001111011111101001010101101110010110000011010011011000100001010101011010001101100001001000000110111001011001000110101100110010010001111101101010101100110111110101010101111111101011101100001000111110000101010111110101001101100000010010001100000100010010001011000111111101101011110000101111001000101100000101000010011111010001001000001101010011010000111100111111101101101110011111010010110011001011111110101010110010100100111011111000000001010110110100011001010111110011010000110010001011011100100011010101101110101001111110001101100100110011100000001001010100111101000000101101000000110010001000000010000000100000110101011100010110101100010111010010100000111111111010111111111110000101101110110101110111001100101000010001100001110110000010110001001111010001110111001111001100001000011000110101110000001100011110011111011110010000010101010010010001110001110110000011110000111000010110011100100101111111110010110101111111111000101101011010010110110010101100011100111000100100001010001001100001001000010011001100001111110111111011001000111110110110010010010100101001100001111001001111100001001011011011101011101000100011000011110101001011001111100011101101000000001101011111010100011111011100001000100111101111111100010001111000100111011010001100001000011110101110011100110100101010001101101001110010101110110000010111111110101100010001001101100101000010110000011100011001101000011001001001000100001000010001100001100101000110010100011110111001101011010100001111111100001100110011011011011010111000100011100011011010010010110101101110100010011100100111000011001001101011100011010111011010100101000110000001100110001011011011001001010111010000001001101100100101100101001011101110100000101001111000001001010001010011110001000100001011100000010110110111011110000101101101110000100011100111110110000011000110010001011001011000001011100111001100110110011001101010001010010110100101000000011001001111010111001100010100100111011111000001000110011111010011101100000010011111111100011011001111001011000100011011100011110001000011101010111110101000010010110100100101110011010111101101000101010111010011100001110111011000010101001101011110111101001110010011111011100101000101011100011000010011100011100110111001111110010100000101011110110001111001010001010011000001000110000110000101011110101111010011001101111111101111101001011011100010111011111111010001011001100111101110001100110101110101111110101110011111110100111001011010111001010110001100101011110000010110100100000011100011011000010110011111110101111000100001001101011001100111001111101011000001010100111100110100010000100000011011000100100011101111011100111011001011100010100111011001111100001010000011010010000010000101011100100110011000010100111001011000100010001001110011010100001101010010011001000110001000101101100001100101100000011110000110101001011100001011110000100100101101001101110100000101100001001001010111010011111011011101000001001000101110101101010000101110101110011000100110111000110000001101100101100110011010100110111010000101100100011101001010110100110000100110111100101000011010010101110001011011101101110110111101011110110011101010110010100111011111100001100101100001111100101011110100110010000101011010000100101100110100101011010010100000011011010111010111101010100011111111000111111110010100110100000000001000000110101000101011110100000111010011101001001101101011111111100111100001100100011011111101001111110110110010001000101111001001111111101110110101000000010111010111001011011001100000001110100000010110001000101111000110111110101001001000110100100010000111010011110000001010110000101000100010011010110101000000011100001111010011010110101010000111100000011010100111001001111111101111111010011010000011100110110111100010111000011011101100100110101010111011100001110100101010110011001011101011010111000011001101011011001111000111011110000000000001000011000100100101100101010101010011110011011011011000111001111101110100100111001111000111100011111001001011010111110011110010010101100011110000101001101001001111101000000110110110010100110110111100110010001100011000001001001101001010010001010100001110110000101001011001001010110001110011011010010111110001111111101011111001111101000110100000100000111010010000100111001100100110101100110001101100100000111111010010011101011111011111100101110011011001001110111011000010111111111011011101110110011110011110110000110000111100001010010101110011101110111011111001101011010010010100001101101111101110100011101001000110100100110000101111010010111101100111110011101001010000101000111010011010111111001101110001010110101010100000100001110111011110110010010001111100001101100101110110111100111110111001100110101100110011010101101010010000100011001010110000111100100001101011010001110101100000110001011000100011001110001101101011100100101000001101111111011000010101000101101101011111001100100010111001000011110101001100000111110110100001001101011011110110111111011110110101010001110001011001101010100001010001100100010110011111001110000110001101010111010101001011010010000011001101111110110011011101000110110111110101011101110101000000010011010111100100000011010000111011111000100111010010011000110000000001100101101001011100010111101101100101010011101001000001001001111100011001110111010010111110111001111101111110100100111011111100110000110000101110111110110101100110010101100000000110100110000010111001011011100111011010000110011010001001010001100100011010111111011001111110110010011100101010111100101001000011101010110010110000111111000011010101000011000111011011000010101110101001001001001101100000000110100000001110101101010001110000000010111000111101100111000011100101111100011100010110000011110101011010010100111001110010110001100110011110101010000111100100101110100110110001010110100001000101011001010101000000111100000010000100000001111101000100010001001110110001111111110111000011110101011010010110111001011011000110111110010011101010100011100100011101001101011011010011000011100011011101100111111101001001111110111100100011001001000110001000111010111110001101111000111111001101010001111111011010011010011110111011100100101011111110111100101001010000011110100111111110001111011101101010010001001100101010000111101111001010110011111101100010101001101000011001101011101010100011101010010110000111101010010011101011100111001000110010110101001000110110000111101011011010010110101001000011001011111100111010011001001111000110001111111001111111111010101010011001101110010011000010000010001101010110111110100001001111100110001100011011111001110000011111000001100010001011110010111101110011010100011101010011111110000101000101101010000100001100001111101111000000110011001100000100011001001101110111111111110110100011011111011101110111110001000001110011100001000001111001101000110001101110111110101110101011100011101010100011000110101111000011100011100111101110111111010101111011001000011101101101001100001111101011111110111010010001000111100100110111101000010100101111100001110010010100001010011010100010101010000010101000111101101110111101011000111101010111001101000101001100101100100110011000010101110011001100010011111100110000001111100101010111110111010010111111010111000010001111001011001000110000010111001111001000110000110000111101101100101000111100000000011010010111000101101000111101101011110110100001000100011010011111000010101001111100001001101001010100011011111110010110110000111110111100011101100111001111000101011010001000110100000101111010111001111011100001001010101000001010101100000011010000110101100000000000110101001011001110000111110011001110001101100000001011000110111111001001001010011111111110111001001111100011010000010101111111011000101000001110101010011101000100100000111011001101011110110111110100101101000100101110111101111100011100101110011000111100101111111010010010001011001011110110011011110010110001101110101110001100010100101000001010000001110110000000000010011111101100001100101001101000110111101111000101010001100101010011100110010000010100110010001000111111101101100101000100111001110111101110001111001100010111101000010010101110110001001101010110110110011101101110100101110001001000111110111011110010100001101000100101101011111001011101011111101101101101101010111011101010111101011100100001101100001110011101111111111101101000100101111110111101011010011111101111100100000101010001111100001111011101000100100011001010001111001100000101010100101001000011001011011010111010101010101111100100000000000000000001111110111000010101001001010010000100001100111010010010011110101001110100011101111100111011110011111010101000110011110100001110001011101111110101010101110100001111011111101110011011110000010010001000011111110011111101100001011010101110001011101110100111011000101001010110111100011010101101110001000011110110001000000010011101100101010101100110101011111011110010001100110000011110000101000100000000011101100110010111011100010011101011101111101000001011100011101001011110110011011111000000011110100111011011101100010011011111010011000101000100101000001101100000100111101110111010001000101010101000111111001010010100010001000100011010100001011001011001011010011010100001100001100101100111101110010010001010111000111100000000010101000011001000011100001101101000001000010100101111111100101000001110011110100000001001010011011010000001011110000001101000010011011010111101001101100000110100101011101010011011100111111010001010100000000001011010100101101100100111010011111010000100010100110101111010100110100000101001111100001101001011111101111001001101010000011011110101010001000001000111000110001111010101011110011011000100101101011010001111101000100110001110010001011100010110001011010111011010011000011100010010100110111011011100110010010000010010111111110100010000100010001101000111001101010101100101001010111001001100110011001010100000100101001001101011011001101010001000001001111101100001010111010010011011011000100010101010010100101100110010011101000010011110011001100011100110110111110100101001011001100011110001111111101100101100111110101110001000011100011110000010111111010110110010000011011111010101101001110001001100010001001101000110100101010101001100101000010001111100110010100111001011000101110100001000011111011100011010110011101101011010011011011111000010111010101010010010011111101001101001000100011001010010011011001100101011110010100000111101010100011000010111111001101111001000010010100111010011101000010101100101111010001101110110010001000001100110110010100010111000111010101011011000001101000101001000100001010101110000101011101100100101101001010001010000101000111001001000000101000001000101111010010110001000000110001010011111100000101100111101110000101010011000011011011001001010011000010101110011111001111010111110101000001101101010111011111101100000010010111111001110000011001010000010011101001000100001100011010011011110010010010100110111111100100001101010101111111111101001111101011010010110010001011110110100010010000110010101110101111010000001111100011110001101110100110100110110010100101011011111110111001011110101010101001110111110110111110110100110000010001111101111000111010111100011100010001010010011100111101011111100011101011110100010100100111001111000111010010001001011011101101111000011110001111100011110000011000101001000100101010000110100000000111001111010010110101111010110101011110011000001001011111001100101010111010001111000010101011111011000000010100101110001000111110010111010100111010010011101111011000101001010111100000001000101000101000101111001010001110101111011111011110100101010110000110101111111010010001100000001011001010101011001001101101110100010111000010001110111110000010010111000100100010001010110110110111101000100100110100110010111100111110000000010000001110000000001111011110000010110111010001000001111101001100110000100101111000001010000001100100110011111001011001000011000110010010111011110010100010111011111010111011110111101111110101101000000001111001101111111100110111101111110111101000101001110111000010111011110010001101010011011000011101100011101101001101111000100010000110010001100011100010011101101110101111001101110010000011000111100100011101101100100010001100000011101110101110100011001010000010010000011100101100110001101100000101001101101100100111000111111001110110101000100011100000001101011010001100000010111100110001011111001010000101001001100111100101010111010010110110011100001100110011001000101101000100011010000011001001101001001011011100111001100110000111001011001100000010100000010001011010110001111111001011000011111110000011000101011000000111110000000110010101000101111111000001011110000101101100111101000111110011100000001100101000100001110000011000101011010110101101001010110010010000101101100000101000110011010101010100000110110010101011110100000011010110111011011110111011001110011011100110111001000001001100101110000011011000111110111001101010011101001101000100110001111000111101010111010001001011010110111001100000111011010100010011011110101001011010000101010010111100101000100111011111111101100111011011010100001100100000000000100011001001100111110101011110001100111100111010010101000111000101111100011000100001000001100010111111101000001010110011110111111001101101001100101111110100000011101101010011001001111101110010110111001110001111100001000010110000011011110011000101001101101111100101001010110000101001101110110001101011010011110101011110010111110000000001110110001111110011101010010100001101111110011001001001000010111001011010101100110010000101101111001001000100110111101011000010001000000111110010011000100100011011000011001100101100100001010100110001011010011111100001111001000100101010001001100111111110001100001100010001010111110101011111001101001000111010001111000010110100101010010101100010000100010000011001110001010111011001111101111111100111111111100110101110111011110100100001010010001011101101001000101010001100101011101101010111111100101001110110010100110100011111111111101110101111000010010011111001110110011110000011010000000100110001110010000010101001101100110011011010001111100101111001010100011111011001000011101011011000011000001000100010110111111101101011011011111111001001101100010100010010101111010100011101001111111011111100110100001000100101110100111001100100111101010011101001101101000001000001101111010110111001001110101001010000001001100110010111010111111000110011001101100111011100011101100001101111110001101010000000001000111100101100110000110111110010000010111100110011011000011001010110000101110110000010000111110001100111000110100110011111111101110001011001000111110101001010000101000110011111001101101010101010101001111010000001001000001110001001011000100010010011001101110110000011010010000101000100101001011010000110101010011010000000110110001010010100001111001101000101001010010001111001100111000100101010011010111010001101110110010101000011001010011010101010100100111111000001001011010010100101100011100000111110010100110000100000111000110111101110101100111101101100100110000011110110100010011101000000100011101001011111101111000011000010001010100001011010010110001111000111001011101110011111000111111100101101110100011100001101001000001100011111100011111000001100101000001101010011011001110110100010100011010011011110011111000101110000111110111010001101100000011010100011111000001011111001111111111101110010101101000001101001110111110111100010101100010010001101110110101100011001111001111001100110011111001110100011110111100111011001100000101010011000111111011000001101011110011101111110100101011110011001111000000010110011110110110000110101001010111100010000100110110001111110100001011010001100010110010010010111000000100110111110000011101011101100101111111100100000000100011011011111000100100110000111000111110101111110110100110001100010111110110100100101101110001011001001001010101010101001111000110000011011000111100101110100101101001111111110111101010101110010101001011100111000011011000100101110101100000011011000011100110001110000111100011100110001110100000110101000011100001010101101111100101000100001011000001111110011011101110101000111001110001011011010110111011011100100110101111101010011101011110010101000000100010110101100110001101001101110011111111000000011100111111001111101101101100110011001000011000000100001101100101001110001101001011011101000101011010010100000100011000111010000101010100000110111111101111111001100011000111100000111100111010000001001110001011001010000111110100100000010101000111100100110011101000110111110101111000101011000001001010001101101110101111101010100101001111000010100000011010010000110011100101110101000000111111000101111010001010111011101011011010001111010011111000111000001011101100001011001100111011000100001001111101110010011001000010001011100010110011100000110100010011110110011000010010110011000100010101101100101010101010000000111101100101111011010001110100101011000100001101000000100001010001010101111100110010101111010100110000001100011011111001010000110100111001110101110011101000001000001000011100111010000000010001111110001110110011001011110010111100010110110111110111000100011101011011011100111110110111001001010011001001000111111000010110000110110000011100111111010010111001100000110111000110101010010100100001110001101101100011110111000100000111011101001011101111011011110100000100001011101101010101001010001110100011111101010001100001110111000101001010100010100111001011110001001111010011001000010000011011010101100111100110101111000011111001111011110101100011001001100010111100011111000011001001001000100000111011001110110110001010011001001000010011000001010000010001111100100110100001001011010000100000001111001010101001111000110110110010010101010111100110001100010110111011110000100101100100111111011101110011010011010111010000000011011010110011111001111101110001001111101111110001101101101111101001110111011101110101011010111110010011101100101001110100110100001101100110110011111101101000010111110100000000010000000011110100111011110000110110001101100001011000000100100001011001111011100001111010101100011111100100101100100011011110001110111100001001101010011101010101110011111010100010010111001100111101000010001010011100101010111101010101000100101110010101010100000011011000000100110110000101011001001111101010000101001000101011000011010101100010010110110101000001101100101110100111110111000100100110101101011000111001111011101111101000001111010111011010010001111101010000110000101010110101100010110101001000001011011001000100110010110110111000011100111011110001111000110101011011000101101010111111010011001111100010111110001100100101010010010110101111111000110110111101110111101001010100101100100101000001111100111110010101110111111100010111101110111111001001110101011000111010101000010011101010111010110011000001111101001111101101111111000011100001100011010011000111010000110101100110001011111101111111011010111000111100000101011111000111001100110100101010000001001111010110000111111010000001101111010101111101100101100001110000010101001010010110011010011010111111000010101110100001001110110001010100000010001011010010011111011101110011011010111011110011011001010111001010011010001001111111010101110101000110100110000010010001001000000111111010101101000100101111011010000000101101000110001100111010001010000110011111111010001111100110000001101101000000111011001101011101110100011101011110000111101110110101110000101100010111110110111101101101111010101101000000011011100000011011001011100001010010110101101101010001000111000001001110110001011101100001100000000110001100111011010010110011001110001101100110010111001010000111101010011000001101101001101000100111001000110100111101001101110110000111000010110111000110011001111010010011110010000111010101010001001000100011100110010000100001011111000001110111010011010100000000000001111011110001011011001011110100101111100111000111010101000000010100110111110101011000000110000000010010100010011101110101110100111010000010001010100010111000011101011101101010000011001001001011100101001011000000001001111110101100000011110010000101000000111100111100111100111110001000110010000011111010010101001101110110001101101011101000000111010000000011000000110100110110001011100110111111110100100100011101011010000101101000110101110110111001011100000001001111011000111011000111100111000100001101001001101011010010111100111111100110111000100111111111000010101010011101101010011011100101111011011000001011000110101111100101100011100101000001101111111001110110111010101101010100100110000111001000110000101001001000111010010000111111111111101010111111001000001101110001011100010011000000000100101000001101001100110001001010000001111110100000011011111001001100110010111100111010100111011111111011110110100101010111001010101000111010101100111101110001011001111110110001000100111111011001100111101101000001001110011111111011000100111010111010101001111000011010100001111101111110010111110110100100011001110001111111110001101011111111101110000011011010001000000011001101001010001101010101100001000000011100000011001001010100011001111110111101000100001101011011000000001010001000100001100001101000100010001000110001011010101011010011001110001111101110011001001000101011001100001001100100110011110000111010000000000010011010101011010101000011100100111001011010111111011001010001110110101111000000000111000000111011110101111000110011000100010110110111111001011011100011001111101101001100111011100000110000101001100001111101001111010000010001010000000010000111000011110001001010001001110100010010001101001100001111100011101110110111101111010100100000111100101111000000111100000001000100000111011001100110011110011100111111101011111110111101011100111010001101101111101000000110001111001110100010101100000010010110011011100111011101001010111001110111011101110100000001000110010000010001000101101010110000110011011101000111111100011110011000010011011100010011010100110010100000011111110010001101000111101110101000100101001110011110100011100111010101100101110100010001000000011111111110010100111000010100110110010000100100011110000110010110001101010111010110000000101101110010111010111110011000001111100101000111110001000100111100011000001100101111001111001010101111011110110011001001000110110011110101100001010111111101001010011001001010001001101110100110100011010110100110110110100101000010011110000010110000001101001100101111000101110001101101001100001101010001000001100000000010100000000110010111101010100001100011011110011000001010011000100100000100000111001101101010110101111001011011000100101011110001110010011000010101101101000011000001111001010100011010010010000001000101010010111010010111110100111110001101101010011101001111101000101010111010100100100100011110011100000000011100111011011111000011110011100000111111110011100001010001111000111000001000101111010011010101011100011010001000111000111100100100111000000001001000111101111010010110110110110110111101100001000110001000000001001011111101111101010011001011001100001100001110010111100001000010100001100010000001100110100011101011000101011000011110110110110010110010101001001000111001110011101110111000010010100101101001101110011111000001110000110010110110101011111100011111100011001011100110110001000101010000001000111100010010010100100110100100010010100110100010001000100111010101000110110101001101001000010000011100010010101101110111111101111101000111111100111011101101011101110010011110100011100101010001001100110010101011011001100000010010000011110110000000100101000011001110110010011110010111101001010011100011110010111111011100110101111111100010001111101000000110001011011110000000110100010101100110010000010100000101110000111011001001001011010001110111100011110000100100111000001000010111111011001011010011100110101010011011001110111011111000100110010101000010110001010100111000101010000111111000101111100111010111111100011111100010100110100000110100110110111111000100110110110000011110010111110000101100111101101111100111100100000111100011010011011000100011000010001101000110101110100100100010111011011011001100110111011100011001101011100001111000000000010100011001001011111011110110111101011011000110111000010110111001110000011110101101100110111110101110010011010000100101111110001001110011010100001100101011101011101110000001111001000001000010110111110110110001100110011001011100010010100110111111011010001010111011111001011011000110010110101101001100001111011011100110000001111011101000010000001101100000101011000000111110011000001001011110110010101110101010100001101010110010101001111100111010110011110110011111101011101010110101111000101111101101111000010011011100000011110100010011001010000100010101001010100010000100010110010100001011101010010011101100001101000111110110100101101001101101110001010110001010111000111101000100010101110011111111000111000000001001001110101000101010010111110100101111010001011101010110000101001011010001011000001111011001011000111110011110111111110010001000000111010000110111101101001111111100100111010011110000101010111100001110010011110111100001100011011111000000010101100000010000010010010111110011001011101101010100110110010000010100000010000111101011001011010000110101101101110000000010001011101010011101010010110100001000110010100010101110111000000010101101101100101101011101111110010110111110011100011000010011100101100001100101011000100101111010000010101010000010101010010011010011011111000011101001011111110001110100101011110111000110101001001010110010000111001101010000010101110011001011011110100011011100011000111011001110001110110110001010110001000111110100110110100010011101010100010100110000001111111011000011101010101011111001110000111011100000111011010111000101110010100111001101101011100111011100111001010111100110011100101010111000100101110001010101111011011100110100001110001001000111010000100011000111101000000000001001110010110100010110110110100101001110001000101000100001101110001010100100101110101010010010100111100001001110111000100000010100101010001111111001101110000010111100110100000000111100011010100000011010010000100110110001100101110111010100110110010010000110010010111011011010100111001010011101100011111001010101011001010011001001001100001101100010100110100101010101010001110010101100000110011010111100111100100011010110111101111011100101000000101100110110100011100100101011011101001000100101010101000000110001100000000010100000011101010110011001111011101101101000101100000110111010010111011110110011001010100111101011010010110111100100000001100110001011101000100011001011110001011000101011110110111010100011111001100000111010010101101110110100000010011100111011010000010111000001101001101101000011101000110001000101111011110011100111111011111101000111110001001100100011000010011001010100001110010111101000011000000100011010111010101110101011101111110111001000110101010111110000100100000000110011101011010000000000000001000011101001000010011011100011100001011110101110010100111010000010010001111100101001110110110010100011011111101100000101111111100101110011110110111000010110010101010100110010110001011111001101010100010001111111101001111001011110111000000100000000010011100010010100111001011001011010101111100100100011010110011001010011010101101101011111110010100101011100001110011001011011110011000000100101111100011111100111011110010000101010100010110100000100111100011000001111100111000111010110001001100011001011111101010001111001101011011000101011110110011000110111010000000111001011110000110011000111101110010001000111110001111001001001000000001011101011011101110100101010001011010011100110001011100000110011101111111001011000111001001010001001000010111011101001001000110101000101011101111011110101111111100110100011000111111101011101001111110010110010101000111010110110010101000111111101100100001100101001001011000111010010110111001110101011010000010101001001011111110010001000010011001101000000001010000010010101010010100001001100100110101101001111010011011101010010100000000000010110010111001101000110001011110101001111101101001101010101111110000011001001001100111011101100111111110011000111010110111110001011110110001011110001011110111111100110101011001100011110001100010000000111111110001111001000111000010000100110001010001111101101000101000001111100011110101001101101000111100010010010110000010110000011111100110100011100101011100110111111111011000101111001110010100011110100001011111011010011100010010000111000001001011101111110101011011101001010010001111110101111101000011011111010010111100010110010010000011010100010001010011110000001001010001000001110010001110011001110111101111011000011010000001111101100111000101101101011001011110111000000010010100110001011011100000001001110111100100101000010110000011110101111010000011001001000101110101010110010101111101001100100000011011110011100000111111100101110111001110110010010100110111110010101011001000100101001000001101001001001011000010110000000010000110111101100101010011011101010010000010100001011110110011101110100000011110000110101000111001111011101101110101100000010100100101111111100110100001100011101001010111110110100111110110001001101100100000110010010101110101101000111000101000100110100100010000110000001110011010000100100001000000001010100011110000110101110010101011000010001110000100110111010011110110111010010110000100010011100000101010000001111111000000001001000011001000011010111000010010010001101001001010011011001001101001110101000100001011111111001111100100101111110101001111000011110010100111000110100101001010000110101001101010001101001110110000110111110111101001001000111011101001001010110111110001110101010001000110110000001000000101101111111001001010000100001011011110001111101001001011000100000001001111110110000010111000111001001101100101000101010011001110111110001101001000100010101001010010110110000111111100100100110110110111111000000010000011110010100111000100011111110010011010100001011101010000000111110010011000010111011001001110001000101101101000101011011011111100001000110111110111000100111111010101000100100100000100000101010011010110100101000010100001011011010101010110010110000001110110000111110000010100100000111000110111101100101101100011010011110101110101001000110111110110000100010111101100111110001101110010011101001111001000011110000001101000111011111101010011010000011111000010010000111000010011011111001011101010100010110100111110111100101101101101011100001101000100101111011101101110110010011001001001111111000001101100111000110100010000000100101111100110111110100010100110110000011111100101010010001000111110110111101000101101011111100011010000111011001000101111011001000110101010011100111101010111111011010001010001111111001100011000011010100000011011001110100100110110101000001000001010101000110010001000110111101111100000111000111110100110111000111000001111110001110001000100000011110111100110111100011011011111100011110000101111000001010111101110001001110000110000000000000100011001100000000101001111000110010110001110010100110111110010100000110111011011000010101111010011101110100110111001001101011001111101000000011011101100101100000011011001001011000010101110011110111011010010011110001100011111000000000110011110110000000000000001001000100111001001010001100010000111111110101011110010111101100010010001011011101111011101010110010001001111001001110011000010010100100100000011001111110010110101110010111010001100011010000110111101101111110100101100011011001100010101011011101111010010001111100100101011001110101100001011000101011010111010101111010010001110100100001011100011101010100010101110010011100001100110000110111100001010100001110110100100010110100011100111010100001010101011000111111010001010110000011111111111101001100001010000011010101101011001010111100010111001001100000101000100011110000111101100100000010101000001011101011111100011010100011010011101100100011000011000011110010111001110010111101101011000100110000001011000011100000000011010000111100101110111000000011000111101110101100000111111011000101100000110101101111001010010101011000001001100010011101101010011101011011010101110111111000110100001110111000110111000101011000010101110000100001011011001000100110001010111011011101111100011010010000100110111011101100101100100111100001101010101010100000110000010111110111111100001001100111011001001001000000101101001001101111100101011001111000001100000110110110101110100010101001101100001101101011010001100010101100001000100010101101111011100101001010011000010001000011000110101010111110110100110100101100010000101111010010011001001110110010011010000111000000001010110100101101011100000110110010101000111011001000101111110001110000110101000010000101000011101111010001001101101011000000000011100100001010011100001100110001100010011001100110101110111111011000110110100011111010110001001111010111001101100010000100110101101001010101101000000001010011000110100011000111111101000101001010111000010100100000010000001101111010101101100101000100100111001001111111101101110110001001100011011101110110000100000101001011001001111000000111101101101111101001011000011000001001110001110111001010000100011010000110101011111001111011110100011111000101111001010100000100011110101110110110101101111001011111001010000100100001111111011111001001011011100000111001010001010001100000101001101000011110010101011010001111010000101100111000011001110110101111001110100010110001001110101001111000010100100111010010011001101011101101100100010111101000001100101011111010101000110111101100011110011101101001111110001111001101000100010011000001010100011111110011000111110010001110001011110001011110110010010110100101011110100101000101000010110000010110110011110011110001100001110001001001001010011001100100101011000100110000011011010100001110100100101010000010001011111100111101010110111100100110100100110110001101010000001101111100011101110101001000111110110111001111100100100101000111111000000000010011000111011110110111000000100110000100100110101011111011110001101111101100001101110111101101001110010000111110010101001110011101000110100000001110100000000101111001101000101010010010011010111111110100101111010110101110000111111101001000101111101011010110000001010110101010110101011010000000001101001100000001011111111001001100001100001101011001110011001111001011111000000010010110100111110111111101001100110001001001010101001000000000001101100001000100000110010111011101011011000001010101011000001111001011111000010001011000010011110100100011001000011111000110110100011000100101000110101000010010111011001001010010110000110001111110101000000101010011101111010000100111111011000101011011000010010000000111111000111100011011001101101011011011001000110111100110100011101100011110101001011111110101100011101001001110000100110010011101111010001111100011100110000111001011000011101110011001100111010010110111101111011010000111010101101000101101011001001000011111100010111101010001111010011110111011010010111100001110100011000011010010001100000001010000011001011110111100001000001111111011101111100110011101000001110101101010011101101011101010101100111101111101011010100010101010110011110000011111110110110111101111111001011010011000101111110011100110111001001011111110000111000011010011010010110010000111010111000101010101011011001010000110010100110001100101101001001000111101100100111011100000111101010011100010101111010011100010100111000110111110010110011110010101010111001111011000100101010101100100100100010111111000110110101110100011000110111010011101101111010101110101011110010111001001010100011100100001011110001101010101011001101100111001000010011001011010110000100000010010011010110111000001000101001011111101111010101100001101110101000100111101100100010110100001101100101100010010101001111011011000110110100110010001110001011011101110111101000010110101111011100111101101101001101010011011010011101110110011111111110000001111000011001000000101010001010100001010101101001001000100110001000111000011011000000011110001001011110000011110000100001101000110110010101000010101011110110111111110100111100110100000001101111010101011110110101110000000011001111010110101111001001110101000111110110011100111011010100110011110111110100100100010101111100100100111110011011111100110110010010011100111101110111101000111011110111100011101111001001000111110011000111001101101000100110001101000011001111101101111000010000111111011000011111011000101100010101100000101011011000101010011100000011111100011101111000001010001000011100110000111011110001111000111001000111001100111011001011111010111110110001101000111010000001100110011100111111001011110111000100101100011010001111010110011111110110010110001000100011100101000010101100011110001110111000110011000011100111010110000111110011010010000001100101110100101100110001011110110111000011001101000000000010011011011111110111011111101011101111111110111111000100100110011010111001001110100100000100000110101100111100111101001010011110001001101110101010011000011101001111110001001010011010001010011011101101010111011111111110101001100001111010001100011000101100101111010011010001010000100001011011000011100110110110010001111110011111011001110011110111001101000001001001110010100101011010011010101101111100100101011100010000001000011110110011111011110100111101110100100110110011001111001111010110010000001011101100101110010111100101110000001010001001111100011010001101101011101000100001110101101000011011010100100000011111001010001101010001001011011000110001111100101111000111010001001111111000101010010000000001010010010011001101100011100110100001100101001001100111111111110010111001110000011000100011000100101110100111111110010100100011100000111110111001011100110000111110001011001101101100111011100010111110011100011000000110000101101101000100001001001010010101111011100111100101100010000111101011000010111011010010001111100111010001110011011011000000101011101100111001111001010000101101111111001101110110001001011101011000011011011010110000001000110100111010001100011100100110010101101011010001010100010011011011001001011010100101001101110110101101100101010000100001010010001010100111010001111101001111110111100110010101111010111101111001110000101010100010001001111101110000101100011110110100111110011111101011100001010111101111100100110000110110100000100001110010000000100000001101101011000001100010110001001101000110001000110001101000011100010001001001011111110010100111110111111111111111011110011111100101110001011111100001101100010010011000111101000010011001101001010101101001100110011100101000000100111110001100100111010011001100111111001001001001000111111110001010101100110011011100000010100100100110111000001011010001101101011010010111110011000001111001111010000011000111011101101011101000001011010111011010010010000010111001101010011110100100111011001100001111011101110111111110010100000101010100011110000011101001111010101110100110000001011010000000101001001111100111111110101101111110110010110101001001011010101011010011110110111000101001111100111101001010011110010100101111100010001001001011000100110001110010001001000000001111000010100111011101000000101100101001111110001110010110011011111011010101010110010011111110101100100000101000111011001110011111111011110001010010000010000110101011001011110011110111000100110110111101101111100010100100101111101011000110010000000010110110010111110001101000010110111101110001001111000101110101011111100010010101101111011101111001100101100001010110011100101000111001011110000111100010100110111111101010110010100100110100010001011110100100111111001110000101100000011110100101111011010110001110101011001000000110001011111110011110110101000011111100000111111101000010111001101111000110110111110001010010000010000100011010000000011011100011110101111011010110001101001100010011001110101101100101110100011011000110000101001010011000010100100000000100010100001000000110010000010000110010011010010101110000101011110000010000101000101001111000010011111010010110100001011101110000011111000111010011110010000000111100010001001000110011100010000100110101011100000100101000011100110001101111101110100001010100011111101101011111100010010110111001110000100010111111101100111111011011100010100100011110111001100001000110101010110101111110000000100111010001000101010110000101111010110001011111111000000110111111000111111110000100100101101011010100111100110010111011001100010100000110011011001000011100001011100100101010101111111101110001000111010111110011000101111100000110111011100111100111010000010011000000010100011111000101011101100011101110110010100001010010101101010001000101101100000111111111111001111011001100100101101100101001100110111000111000100010011010100000001001000011011000111000100001100000011010101001100000111100101001000111010110011110001100100001101000000110010011011001001010100010000001111100010100111111010011101110001011011110101011110111111111100101111110101100101101110110011010001001000101101100001100100101010101011010111111000000010001010111111101000100111100010100000000001010101100100101001000110110111010011001101100001110111001101011000110111111011111100110100011111110001100111010001010000000110101111100011100011001010001001011100010100100100101001010000111011010001111111011101111110111010000011101010010011011111011010101010100011010110011001001010011000110010001110100000111001110001101010100010101001001100011000110100000101110001010111101010111010010101011000010000000011111100010010101111110010100000111100011011001110111001011000110100111001011101111101100100110000101000111001110000001001110110110001111101001111100111110001111111101001001001110110000001101010000111010111000100011111111010111011001110110101101111011100110101111011101001111111111101000001101010001001100010111100000010111101100111000111000110100010011110001100011101101011010110001001001100011100100010000000110111110011001100001001111011000111100111100100011111110101000111010010001000011001010001111010000101111000101011101010101100111110111011100010010000100000001110111111011011001000010000010101011001110010000111010111000001001110010011101110011000110100101000010011110111011011101001100111101011001110000011001111001001010110010011110011010001011010101010000100000000110101111101000110100000000011100101010101111110111111101101000110010110111111110101000110010000111011101010000101010110010111111000001000010100000010110110010000000111110010100111000001000100000000010000001001001000100111111001110100010110000111010011000111110110010010010001110000110110011101000111011011011011000000010111011011010011111100000011011000000101110000010110101111010010100101010100010101110101010111000011001000001011010010011101100100101110101011010000001101110110111011001011100001001011000101100010100001010000011001011110010111010001101011001110100110001101001100001001000101011000111111011001110011101110010100100000110010111001110110101010011101000010100010010101011110001011100001111110111101011101111001011100010110101111101000001001111000101010111000000000100100001011110110110110010101011000001001001010010011100000101110110101001010111000110110011101011110101101010011100111011100101001010100100100011100111101111101001001111011111000000000010100101010000111111111000011010100111101111101101111000111010111111011011101001010001011111101001101111110101100011011100000100000100111000111110010110010010001000000100000001101001010110110111010011101110001001100010001011101000011000011110101111001011100111010111001110000001000110001101011100010110110101011000110000110001100011000100001101010011011101100011000000010100011110000011111101101011010101000100111010100100010111101101010110001010010101100000100011011101100010101011010100111011101010110101110000100000101000010011000101001000000001100001101000001110111111000111110011101000011110000011110100010010111110010000111110110010000011111000011101110101110001110010101111100000101001111101001100110001111101001111000010010101111110110000010010010001111010010101001111010001000000001100000110011000110101100111011010011010001111010101001001011100111001110111000101100001010101011110111110010110101111001010101110101010110100000001001100101101011100001011101110000010110000100111101000001000000000100101111001110010010100000000110001000001001001101110000100010000010100000011010101101011110101100000110110110001001001111111011101110110001100001001001001000011000001110010110110111001000110110111011000101100110001110011010101101100010110000011010110101001100110001001001000101010100001010011010000110101001101000110001001001100110000001001101100000110110001000010011111101001011001001000101010101110101001011100011000010000100000101101101111010001101011110000000011010001000000111010011111011101110110111000111011100110010011010011011101100111100111111010001100001011010011010111111010110111101110000111010101110010010111101101000100111000111101111010101110111111000110101101111011010110100001110111001110001111011101111111101100111101001100001100000001110100010010110000101100000011011000111001111100101000110101011111101011010111001100010001011101101101001100110010111111010010001110010111010110111011011100100010011000110011110100000110100110000110001011100100100001000011110000001111000001000001010010110010110110011101000000100111100110101001011001011111111000001010001101000111101000011011110101111100111001011101100111110101011101110000011111111100111110010110111001010100101011101001010110010101001001100110001110010001011001011000010111100001000010110111101100010101010101011000000111011101010100101000101100100011101011011111100001010111111111111100001001101100111111101001110100101110001010110100101110000111101000011001000000111100111010010111000001110111111100100010000101011010100101011110101001011000000100011010101101010001101011000101110000001010011010101111111000010101000110011001001110001011101100000011110100110100101001111100110011110010001100101011100001000111011101010111101011011011011101101011100101001010101110110100001010011011110011001010010100110010101111110111111100110100000001100001001111111100111000100101010001011000110000000001010010100001110011001111100101000100011110110011100011100100011011011010010101110110111111010110111011110010111101101111011111010101110100111010010101100110011000000001111101000001000010100100110001001110001101011001001101000000101001110101001100001001111010011110000010111010111101010110100010100111101000100100000110001100111110101110100001001110001101101001101001100111000000011101111011111000011010001011001110110110001011100000011111110100101010110000101000101011001101111110000100111110011111010011100101000001100010000101010100001100001111100110000110101001010001101110110101110101101110001011101111101001001010110100011110010110000100011000101111011011000101000001000101011110010101110110111010011010000110000100110100100011011111100110100011111100101111000000101111101000111011011001110110110011101100001110110100001001010111111000010001000011101000000110000000001000000111011010110011011111110101000000000100011100001010100111100011010011010111111110101011000000000010011000000111110100111101011110010000001100001110100010000011010011110000101000001111100101111011000010000011111101010001100100010111010101001111101111000100101011110010011010100101011100111101011111001100100000101001110101001110010010001001100101000101001101101111101001011011010001100110100011100100000100000110101110100000011010111101110111110101010000010001110000010011100010101100101110111111001001111100001100101001011000000011111111111011010010010010100111100000110101101101001000001100000101101011111110000100100010011011011110110111000101010100101111110101101111110010011111000111010010110100110011000100001110011001010001000110100100000000111110110000110010100100010001101000111110001011111011011111100011110101100100000001100010110100101010010100101110111101110011100010111110100000110100110110010111111110010101100000001000001010010101010101000111011110110110010111100011110101100111001111101010101010010000111001011101001001011101111011010001100101110001110101101000010111001110110111100010101101111001010010010000011000001000111000001101111101100111001111000011111000110010001110010001001010011110111110111010010111000110011000000110101000000000100010110001001010110111110001101000011100001100110011100010100111000011111100101100101011001101011110100010111100101110111101000011111011000010111001001001011000110100111101011000110011101111001011111111010100101100110010100110111100011000011000110011101011010011100101110111010100001100110011000011101010100011010101101100111101010001011001001100110110011000011111000111111110001100101011001110010111101111100100101011100011110011111100101011010001111001010010110101110001101111001101111011100100111101111010011011001110111101110101100111100110011010101110101001011110100101110100110001001011101111110010001011011101100001010000000100100000110110100001100110000111101101001110001010101001000110010000000110101111001110101010001100101000000101110001010010010001110110010011101010000101110000010110111101010100111111110011001110110000100000110110011100101101100100100010010101000110100000101000000000111101000100111001101001011111100100100000011101011010000000100111000010111010000001110001100011111110111111010111101110001100111001001111111110011101110100010100101101000110100111010010100101011010011101110010100111001111011100101011111100001110111001010111110000110001001101110001010001100010001111110100101000011100000001010000010000011101100001100111110000001111100110111100000110011011001100110110010001000011110011000101101110011000101111100001010001011100111000110101011011000000110111100111000111000011011001101111001101101101110011011100011010100111000001111101100100111010011001100100011001000101110001001110001110001101100000001111000001101011000110011000111101010111011110010011100100010010000000010100011111111111011111111100001110000010010111110011010011111000111100010101111000110101001110110010111111001110110110000010001111010001010101110110000101000011111001110110100111010110000000110101111001110011001011001011111010010111011100000011110110111010000100010011000100000111000110011011100000110001110110111011000101000110110111101101100111000000001001011110100100110110000010010110101100010011111111110111001100010111111001010101100010110001000001011110101111010000001101100010011010101011101110110111011101100011001101000110001110100110100110001001011011101110001011100101111011010100101000000001010000001011111110110010101100110111101001001001010011000111100100101000111001010001101110000110011010100011010110110001010111001001010011100111101011110111001100000110000010010111010001111011111011001001011000111010111011111101010101000011101110001011010110100101110011101100001011100111100100110100111000011001000011101001101001001110110000101000100010111100001101010110110011010001110100010011101010110100001011001100110010111111111000001011011111000001001110101000000011000100001010011111100001000011100000101001001010101011100110011101001100100111010001100010000011001101010010101101111011000010001010001011001100010100110011011000011011111010110100010101100110111011010101000101010010111010000000001011010110000101111110100101110011011011010001101010101011011101100101011100101100000011011100101001101010001010011001111011101000001100010001100101011111000001001111111111010011111100101101011010001100100001101100000111010111110001010100011100001111111011011010010100001000001001001111001101000000101110000010010010000110011100011111101101011010101111000001110101111100000101011010100101110101100000010011101111111110111011100111100000100101111101011101100111011001000011111000011001001100000000101000011001101011001110111110001011110001010100000111011001011011101001000010010000110110010010010001110111110101111110010101111111100011010001000111101101000101111001011100001001011011001101010100011111100001010101001111100000011011101001011100111000001000011110000111011001001011100001101010101011000000110000100000011101011000101111001000101001101100010011111111000110101111001011100010100000101011011001110111111011000000110001011111101010101001011011001011111110110110000000000110100010111100011101100110110001100101011101001011010010110001001110010000110011001110110011000100111011001001111110100001000111000101100110111010011011110011011001000010111011110010011000111010101010110110000101101010111100000111000010001000101111011110001011001110110010111111011111001000111001011000001101010111100010001110000001101010100100011001111111011110011101100001001001001010110001010000101011110111001101101001010000100010001010011001001100100100111111110111100101010001110101111011101101001111100001111110010110101000100010010101000100001011100111110011100000000001011010011010111000100010110011000010111111000010101011110011010011000111111010011100010110011110000010011111110111010100110101111110110011011100100101100100001110101001101001100101000101011111010010100000000110110100111101011110001111110001011011000111001001100000011100010101101111001100110000111001110110000110011100000011001000011011010011000011000100000111101100100101001100010000101110010010010011000100110011101101011111110110011011001101000001110011010000101000000110001101111111100110101000111110011111011110000010010111100000111101011001111100000100110111100111001111101000011011011000100001010000110010111100010111100110101011110101000001100110101011100010101011011000110111010111111100011011100001000001110001101100100100111010000100000010000100011011111110111111111010000110110001100101110011110101000100010010100001011011100101000100101011101110000010110011110101111110100111101101111110100110111010110111100001000000110001101110010011101100111110111010000001100100101100100110101111000010001111010101111111010010001010000100110010010110101110000101000000000000101101001010101110001110001010111000111000000101001110100100100111011010001000001111100001001010111010110000001111011101100001001011111001111111001100011010000111111001111000001000111111110001101010011111001101110010010001010011100101101111001011000001010000011100010001000111100011001010110010010111101010101001011100010011010111111111111011110101010011101010010001011000000011110100111100011100000000100110110001100110011100001010011111001111101010111110111101111100110001100001010000100101010011001110000100100011000100010111110110101000111111000000110100010100110101100110010000100101011110000110111111001110011101010011000010101000110000000110101110011111111110000010011011010111110000110110001111010110111101001000101011001101011110100100001101110101000001001000101110101100101110011001001000001100001100011111000111101010110000011100011111110101010001000011001001011011011110111100100001011111101000111000010101101111110010010010010010010100001001010101000010100110110101000100101011001101010011011010011101101000000010110010100010000100011110001010010011010110111010010110101010101100111101111100100010100000111111110010101000110011110101011011111110111010011010011000100101100000111111100011100011010111000111001100000000110111010111000001010011001011010100011010010000010000001011000011101101101110111001011101111010110011111101000101001011100111000000011101101110110101000001101111110100101011010111111111001100010100101010111010111111101010110100100111100110101011001011110001111000110001011111010001111000101110110101001111000101000101111101101000101001100101011101010111000011000110011100101000100011001101010010101010101111001100110110111111010001100000110100101100000111111101101111101000011110010110001010010111101001110010010100000011011111100100011000111000101000011001001010111001110110000001001100100011001111010001111101011101010010000000110100110111010111010100001111001010101100101100001100001001110001100011100101011001101111101011000001001010011000111011101011100001011000010111111100111100110001101110101111000010100111010101110100010110010111110001011010111010010011000011001011010011110111000000011010111110000110000111001000110111111010000110100111111110110010111000101111111100111111111101110111100111011010110111011011111001001000000000000110110110010001100000101110000000110110011111000011011100100111011111100111110111101110110000001000000100110110011111101011010100001000000101010110101010000001010110100011011001011001011101110000101010100111101010001100111101101100000010100111111101011101100000110110100000010111010010111010100001101010110010001011110000110100101111101001010000111010011110111110101011000110101100100100111001001000100001000111011011011111100111101010001011000010101010101001110110000101000000101110000111011110010011110010100100101101011111000111110011000101010111111001010011101001101011001110001010101010000010111100000000110011110111111011011000100011001000011110011101111101110101110011000110011101100001000111010111010111101011100010010000110001100001100011001110000001000110000101111110000010010011001001111010001111000010110101100110000010111001000000011011101110000101010100001000001010011000011110010111100100000011000010101100000110110011111000000001110001101001001100101111101111100000010110010111111111110111100000011010111000011001010011110101111011001100000000010110111100000110000101101100011011011100110110110101011001111011010010000111010111100001101000100100111100010011011110011111011000001101011110110011000100111101110000000110001000110000110001110111010110000000010000100010001101010011010110000010101000010100101110010111001001110111001001001001111011111000010010000100101010000110101100000111111011110101000000101110101100010110001000111010100000101000101010100000000110100111011101101001111010010010111110110111100110111110100011001010110100001110000111100100101100010111101001101000001000110010100101101110010011001101000101000001111010000000111101100000011100100101011011111000011011111001111111110111100011111110000101100100100110110010101011011111000101010101100110101010110111100011110010101001100111010101001100110101010010110101010101001111011101011000001110001001000111110101001001011101101010011010100010000110010110000000001110000000000000100111000011101111011100010100001111110110110111001011001100000001110111010111011111000110010110111011001111110100111101101100110100001111110001001010101111000001011010101011010000111101101100110111101100100100000110011110101111001110100010010101101110001011010010100001100100101111101100000101010111100001011111101100110011111010110000101100001101101011111100110000001001100101010100000110010010110100111111001010011001000101111001000100000100000111000100110101001001110101110111011011110111110101011000001000110011010011101110010001011010000010111011011100001110100110001111010011010110101101101110000100001100100111001101001010110001101111011011000010011011101000001010011011110001001000000111100110001101111000110011111101000101110000010111001001110011101000010010111100010111001000011101000101111001100011110100011010111111010111010000111001011001111010000101110001110011011111010100001011011100011100101111011110111000100111000010111011010011100001011100100101000011010100100111111111100110010001111111000111110001011101010001000100010111010011010110110010010011110000110000010100011000110011100000000101111110101110010000011111000000000111011110110101001110111100011111100111000010100001100110000001101111000101100000111011000100001110111001011110010000100100010111110010001011001000000111010110000101000000000010001101100000001100011101000001111101101001110011000110100100101011110101101100111111101101101101101100001000111101101111101011110100110110000010011100100010100001101011011010101011110100111101110001111011100001001101000001111101111001110111111100011011010001101101011111100000100000001100101110101100011110111011011101101110101100110111011100101100000111010110110101010000111010011111111010000101110000010000001101100011001011110011100101001101111101111000111001011010101000011101011111001001111100110111110111011110100100001000110000111000100000111011100111101010100111001001111010010010100010111001001011010010101010111101101101110111000110111101000010010110111000110101110010111111110111101001000101000000001100100111101100010110011110111000110011000100110001101111010110111100101000011000000010000101111011100011111001011101000100110011000011111110111110000010111010100001101101110111111111101110010101011000101000000111011011000000011100111110011000110100010100010111111110001010011001000100111010111011001110101100100100100011101010011101100101111011111011100100011000010100001011010011011010110111100000101101100000011011101101000010101000110010110010010000100100000010011001100111100010001001111001101010010111011111111100011100010000101111101001001101100111100101111111100100101001001101001001111010011110101001011001110100000101010001010000001110110011010100110110001110001000011010001110101010011001011111100101001111011101111010000101101010001001100000001100111100010111100101110110111000000100011011110000110111001001110001011001011001010110110001110110011000100010011011000101000111101001000000110111000100001000100011101100000110011011000101101101001001000111001110111001011011101100111110100101100111001110111111011001011010100000011011110111110001110010010100010011101010111100001001011101000010101010010110010100101001111011110010000101111000011111111000110100011010110000111110011000110011101111100011111000010010100000011110000111100011100001100111101011111011110010010010001001101100010001101111011011010111110000101101111110111000000101101101010000001110001101110000111010000110100101101011111110100100011110111100000010000111010100101001011010111010011000010000000111001011001011111000000010000000110001101010000101101001110000110000001111110101001111111100111110010011001110100101001100101000001010100111110110011000110011010101100011011101111000100110111111001011001110001111011111111101101100011111001110011011000111000010010110110011001101001100000101110010111110111010011101010100110110000101100001100111110110011001010110001001011101001100110101111000011111001100011101100111111100011001100011100110110101000011001001001101000001101110000011110011010010000011001001001111001011010011000001101001001001011110111100110101011001110010010001011111111000101111010101100000100100011010111100011101000100110100000111000111011101100100110101000000111100100100101111110000011101001000101001001011000001011101100100001001110011000100001000100011001111110010111011111111011011111101100011101110000000000110111101101111110110111011010111100101000111001010011000110011101010001011101001000100000010100110100001010110001111010011011001000110011100101101010010100110010100110100101110011101011011000100110111001100100110101100111010110000111001000110001100011100011000000000111110100111010111100011101110010000100000001011011010101001100101011111000001111111101000010111101101010011010000011010100100101101100011011100111011100000011110110011111010111000111010101001100000100000010000001000000001110100010011010110110101000000110111111011101110100100101010101001111000001111101000000101111101011100011111011100011111111101101011011111010110000111101111101111001111000110011010101111100110011110010000000011100100110010010110111100011000000001101111101110011101010001111000111100100111100110011101011011011101111110011000100111101000000100000110111100100110000001011001001001001000001110111100010111100011101101101110111010110111110100111000110110100111101111001001111001001101010101111000001101111000101010101110110110010101011001100110100101100101011111000111001011100001101100000010110000110000011000000111011000010001110111000100011101001111111011011111100010111101100010110010110011101001000111000011100010111001110010101011101100010111011010101110111010101010110001111011100011111101110101110100110000010000011100100010011010110100011000110100001101101010101001001000111011101011001011010101000011110111110100111011011011010010010101000010101100000011111101001001111110000101010100100010101110011110110010110001101000100001110000111010101111101101100010101001000010001011101010111000100011000010110001000100001001101010111010100011000100001010010010000011110100111001101111101011011101100011111000011110110110111100111101110110101000110011111110011110011000011011010100101100010001111101001110000001101001001101111100110101100110110010110111011111101100111010101001011001001111101011010111110000010101111010011001001001010111011001010000100000001100010100111001100110110110110111001111110011010100110011010001101001111101011110111111110101100110001111001111000111000100001010011010011110101011111111011111010011100101111011001001011100000101110101010001100100110101111000001101111110111001000101010001000101011000001110110110111100100100110001011110000000001110100101001111110100011100101101000010000101011001000000001000100010011110011110011010111011110110111111001001000100011010101110000000001010011100100000000001010000110100111101111011010010111000001101001000011110101110010111001100000011010001000101111100110010001100011001100001101101001001100111000101111010101110010110101110011011110010100001000111011110101111110011011000010011010000110000111000110101111111000011101011011110110100011101110010100101000001010110001101111011011100001100110010010001000001101010011011110110010010101111000111111011000000111011101110101011001010101011110011000001001011100100011001011111000001000110101100000110011000001011010111101010101111010010110010011010010101111110010100100011001011011010111010101111010011010110010111000011001100010110100101100101110101110100101000101010000011100011011001100010100001100100000010001110000000010100111001000110010101101111000001001111000100101101011010101100100010100000001011110101111101100110010000010101101010011011110111110110111001000100111110010011001101101110101000010010111011010100101000000111010100110010000001000010110010000111011110100100110110000000101110101101011110100000010101111101000001000010011000010011101100101101110111100100000110010001001100001011111100000110010110110010111101100110011110010101001100111101101111001000110000000100011111011010001000001010101100111111000110100000101000010100100010101101000110111110110001001001000011000000010101011101111010101100110011011001111110101111111111101011110010010110111101111100011111100011010001110010111100110011111011010110011111110011010001111010011011101111001011110011010111010111001001100001100100100001000111000100011110111110110101000111100010001100111111010001010100101000000011101000001010000000011010011100001001001011000100011111000001111111010101100110100100001100001111010111111000110111011000111111101101010000001111000001111010000010100100100101001100110000101010010000111111001100100001101000110000111011000001100101101000111100000000101000111010001011110001111001111111111110001111001100000100101111010100011111111010101101011101000010100110111100011100010001001001011110110101100101001011100011101110110011011001111110000000000000101101001000000101000110001111100001010010110110100100001000100011011001011110000011000000011110001010100000011011010101100101001000010000010110010010011111101101110101001111010000000100100100111110011000011010001010000001010000111010000001001000111000111001101001100010000000111000110110010111000000000110010000110110000001101011000100100011000000010111101011011111011101000111100000111111011011100000000101000010101111101001100110101010101010110110110000111010100110100000001001111001110010000100001100101111111111011000010011110111011010000010101011000111111001000101111100100111110110011011110100111010110101101110011101011000011101011100101010011011110011111001011010000000110110110101100111011100110010010100111101100010110100101101000000110101101100110001000011111011000111010101001011000101000110100111011000111011011001001001011100011111000011110100000110101101011111000010101111111110111000001111000011101110011100101000010001011100100001011100010101101001100101001111011000001011001100001010111001000011101110101011100111100001010101110110001101111011110100001100010011011111110111000110101101011100001110110101111100101011100001101101001010100010101011101010110111001000011001100001000111000111101110001100101101011000000101100011011001111001000010000000010101010101001100011010100101011001100011101000101110000111000110010111110011000011101011100001010000111100011000100111111011011010001111001100110011100001000011110111011011111111000000100111010101010001101110010001111110100011001001111100110001001000111000000001010001011010110100000100010010011101101011011011000001110110110101000111010010000000010101001101001111111011000110001000011000001110100101011011100110111001110001101100000011100010110010000010111111110110010011011111011001001111110010101001110111111000011101011110011111011011101111111101010111101111111010011001011010110101100001110011111001001111101110101010011001101101000101100101111100100101000001101000000011100011101101110001011011011001100011011011100110010101100000110001011010110001100101110111000010110100011000100110000111100111011100101010111011001010101101000001010101011111101101110001011000001001101111001001100101000000110101001001011001100011011010001111111100001010111111110010000000000100101101000111100000110001000010010101111110100100110100111100000010010110010001110011111110011110101111001011000001000110100100110001110101011000101111101100001000100101001100000001100001111100000001001101001111101111001110010101011101010011110010111000001011000011111101101111101000111001000101100011100110011011010001000010101000101111010011001001000110101101111001011101001011001111101101011000011000111100110100011010011111100001111011011001111010010000110111001000100001001001101110100111011111100000100011101000001001001001011110110111011011011001110001101110111110010011001010100110110011000110010101011000110001101101111000000010011111000000110010010111111111110011011110011011010111010100100100001010111100011000001100101001110110100101001001011101010011001110001101000101110111000110100011100011100010001000110010110111111101011010101011000011000110111111001010101011110101000011111101010110010100010010101110101100000010101111110001010110111110111000110000110110101111110000111001101111000100010111100101000001110011011000011110110110010111010000011111100111111100101001101011000011010000110011110111111110110011000000010110011111001011001101001010011001111100110111110110101101001001111101111000101110011010000111011001100001011001110111111111110010011010100011010100001101010110001110100110111001011011000000000101010111001010010001011101101011100110101010000000110000011111111010000000101110111000011010010100111011110010000010110011101111111111010001010011100110111100010111100000100000001000011100111000010000000100111000100010111101010000001101010100111101100011100011111011100010000100001011101110100100101011101111111000001101101010111001100111110101010100010111010101111010001100101100001001010011010000000000110010100101110101010101100100000110100001000111101010000100110000010001010101111110001011010000010011100110101011110011010111011000101110001110000011101101111101000011110111001110111010001001111010001110010010100100001011100100010010110010100101010101111110110011000110101001100111110110110111111000000100000111011111101100001100110011100110100101101011001011101011111111100001100111010010001101101101111110000101000101011010100011010110011110110110001111011001000110000000111000000010111000010110100010001011011101101011101011011111100101100011011111110010101010000111101001111110000111000110011000100000100010100011100001001011101011100001001101001010101100101010101100000101110000100001010110011110010001110100001001101111001001111011011010011101000100010110010100001011110111010100010100101011001101000000010010000001000110011101001000101011000010011010011000001110010101001011111111001111011101000100100010100110101111100010101101001011111010111100111000011110111101000101100110101001110010000101110101011111001010001101010111010001110011101011101101011000101010111011100011110100100111001101111000110101000101010111100001001101010010101100111011111110101101001011111001000110101101111011000100001101000101010000101010100001100001111010000011000011010011100111001010011001011001011100000101011011100010101101111001010101101110100001101010111000110011100101010100000001000110111001110001011111011100101110111000000010110101100111100010011010111110000000000110110001100110011001000101011001100011100111000100000100110010100001101001110010000111010011100000101110010100000011101111110011011111011011101100111000101100011110010001110001101010011001110011111111001000010100001010100010011011000111100000111001111100010001100110110010110100110010001000100000100010001101101000111010010011100010001111101000101001001010011111110110010100010011110000101011110001000010000001011000111000010110011101011101100100101100111010111001100111101000101101100101010011001011100111100101101101111011011101101100101110101110100110011000011010100010011110001000000100111111110001000110101000001010001100100111100111001101001111101010110000101001100001100011010000011100101100111110000111100010011111011011101010101111011100110110011010000110111110010111101101101011001011010111001110111011100000100011001101101010111100001101100100001001001111010111111000000101110100001110111000101101000101111000001101100101110001001001010111111100000011100100101011111001111101010111101011011001011100001011010011101011000100110110111111000110010110111000111101001110000010000111000100111010110011010110011101010011010011101111001001010110010011111000111101101011110111000101100101000010010010011101001011111101000010111110110101100111010011001101101000100000110111111011101001011001101101111110101110111110001001110011010011000001110111000001100000101100010010110110101110001000000010010001001000000111101100100100110111111101011001111010100000101011001100110111101010010001010001100000001101011001111100110101010110011010011100000110101010010010001101110111110000001110100101101000001101001100100000110001110010001000110100000010001101101010001111111011100111111000110000100111000110100111011101010100010100111100110101111101101100010000010100011111001011011000001101010101100110110011000001101010001101110111111101111001111101011111110000101110110100001110011100011000011001001101001101000010011010001010100011101101100100110000010110110101100001001010011001110001101010000011000100110000000011010000001110100001011111100000010111100111001010001000110001100011000101101101101100100110100100011001110010111000010101000101010000110110010111111101000000010101111110001101001100000000100000100011100011110101001010010110111011101111010110110110011111111011110100010101011100101101010101000010110101111010011101110101111001100001110001101000100000110001101100011111001110000101101110010001000001100101010101111111000001001110011101110001000100000011011010111101111101000010111001110011100001011011010000001001000101011001100001011110101000011011100100011010100010110110000101110010011000001111110011011000100001100111100101000011100001110100110101110011100001101110001001000101100101001001000001001110001111000111001001100110110010000000111110000111010001111101000010101110000011100100011101010100011011000000111100001000000110000000011000001001101010101101100110001000110000000110100001101001111000111101101111000010011111010110111110101000101001110010101010111010011100000010011100111000001011001010001001101010011101001001001011101110100111000100001110010110111000101101010100011100101101110100010001000100110000000110101000011100001110000110110100100011110011011111111001000100011001110001111000010100011010101110111100000011000101001011001100100100001010100010010100111110100010110000101111001100110100010101010100001011000010010000100001111011100110111110110001001011101100111000010101110100000101100111101001011101111011001110111011110000010101010101011111110100001101011110010011000100000011110110000010011101010110011111001101110110110111000010010100010001110110011000111110100001101100101110001110011111111110000100110111111100101011111010001000111110010100111001010101011000110110011110000101101110101111111001101100000010110001000010101111101100110011011001000100100110101101010111101001011100010000100101001100000111101010011100011101110001101111010100100011100001001101000001010101101111110100000000110000011001101011111101001110010011000000101101110001000111110001101101011011101100011011010011001101110101111110001101101000010011011100101011011101110011011100000000010011110001010100001100011011000100010011101010101100110110101111111000011101100000110100100110111010011010101010110110110111010100010111011111110001111100101000110001110100111010100010101011001110110011101010100011001000001111111010101011010110000110110000101010001110101110100001010011110001110110000010111000010001101110111110000001101000010100010101101110101001111110100001110110100010010000000100001101000110010010001001111001001111011110001000111100010001101110000110010011001101110111001011110011001100111001100110000111000111011001000011010100101101110001010111010000001110111011010011110010011000001011001111111110011010100101001100101101111000001011110110111111010110110001011000010001001010101100010011111110011110000011001110010001001000100001101100110100100100011101100100110011100100111111000011111110010000110001101101110010000000001001111111111110000100110000011010111101000111111100010101110110000001110110100010000010010100011111100011010000111110010101110001100111101110111100100001110111000000101100010111110101100001111011010011100000001111001110101101000010100101100100001101100000100111001111011110010101111110111111011110010010011010001111001110111010010010011011111111111000111000111100001110000011010110101010110100001110001000110010011100101000001100111011111111101011110100101000101001101100001001111100111010110101101010010100111110111001110110110101000110010011011110000100011111011011010110111101111011000100100001110010111111010011011010010111011010011111101101110101111000101101110111001001111001011100100100101111000110101010111011110101011101001111111111000010011111110001100011001010001011111011000010001101110001100111010110110101010001101111010010010010001100011011011100110100000001100110010101111001000010101000110011001100101010000100111111110111111011010011010011110100011011100110011010110101001111111110000100111101000101110001100101100000000011010011100111101010001100110100110101111100000100001010111101111011100110101110100001101100000011101010000001001010011001101110000001000010111000110011100100110000011000101101000100011110000010110000100101100111000010010010010001011111010000000101110101001011100110100111011111111001110010011100100110100101101110101111001101100100110101001110100000001010111100111111111011011111100000111001110100011010100001000111000101000100010001101010101110010110101100101001001100101010000111111100110001100101100010011100010000001101010010101101110101001101101110100000101111111111010010010101101100001010000000101111110010001111110010010010011001010110001110010100011110011100100010000111101010000010101010000111111110011110111110100000010010101001001110100001000010111000100010011101010100111100100010000101111100011010110111101100001111100001001110100101111111111011110011101001011101101001001110111110101111100111011110110001001111110001111110111001111110000010000001001100011101001010010111001001000010110110001101100010010101000000000100010101110000111101010000001111100111000110011111101011111100000100101011110010001011111011011011100101011110110001101101000010010000011000100101000111100010011011010010001100010110011100111111010010000100101101111001111001011010101111100111001001010000011101111111101100111000011010111000011000010011011000001111110010010101000000011011001001001001010100011001011101011000111010010000011001111101010000101110111101010101001100101000110010110010010000110011010111111001111000010010110101101111000010010010001101111111101101000011001000011100101101101011111011010111010000111100011001111100010110000010010111100101000010011010111111111011001010000000100110111111110001101111001011011000111011011111100001010110001101001011101000010100111010010001011010011000011110010000100100010000000100001111110001111010101011001001011000100010000001101101110100100011110111010010101001010000001110000110010001011000100101001100101101000000110110010110001011000111111100100101101100010110000110001111110011010100110011111011101100100000010100000110001111000001100100101111110100001011011001110010111001100001110011111100010110101001011001111101111111011110110000011100010011010100110110110110010111110001110000100110001001110011011000100110010110100100011010110101100010110001001100011101011001101101011001011010000011001010100010010001101011110010010001011111111100000000000010001001101101000000111100001111000000110001001100001100010001010110110000100101010011111000001111011101010000110011010110001000111101001010100101110011001011000011110001101100000000010101001010010000011001000101101000011001110100110100111110111111001101001000111111011000110000111011101111110011010101010101101100101101111011001110101101100010000111010011111000110110101011011110010011100100011000100110011101100111010110100001110011000010011101010001011110000110110101111100000100001001001111001111110001110011001101000101011101001010100111000111110110000001001101010110100111001110110101100010100000111101001011001101101101110101110011010110011100010010001111011111010101011110001001100111000000100001011011010100011010011010011011100000010110111101101000101100000101011101111110000001000000111000101000111000001011101010111000101000011001010111001110010111101100010010110000010000011000111100000001101011001100000000001110010001011001010111000000000010110000000110011000110101101111110010100100100000010011010111011001000100000111010001111010001101000010000111011110111100011011110000101011110011111011000111110011110001010011110101001100101011111011111000001010001110010010000101111100100001101110100000010011010001100101101000001110110010010101011110111010110010111000111100010000111010001011111100010010011010001100100100100111000010100000000110110110110110000001101000011000111001011111100001111111101110110101101001110111111011101100111101111001000011111000010000101001011110110000110011101000110000001101111010110011011101011111000011010000100100010111101100111111001111001100001001001011001001011111001110111001110110101100010111101010110110101010000000000000111100001100010111010001010111000000011111111000111011110011111101010001011001101000100000101011110110011110010110010100111100010101000010101000000110111011011000010011110001001010101101110101000011100111001010010000001000000010101001010001111001001010111001100101011011110100110000001110111110111111110110100101111010101100011101011011000000110101101000011100001100100110110011111011101110111000001011011011111011100110110000111000111110101011011111001011100110000110111001001100101011011101100011100001011100011010111110011110101011010001110100110110011111011010000110010100000110000000100011001100000010100000110101111111101100100011000000001011101100111011000101111101010001001101000101001001111001000001010010001010010101101111101001110100011010100110010000000111000000101010100011110101000000110101000100111101110010101000001010010000100100110001100011010101000000100101001101110110011011101111001000110110000010100110101101011111010000101011000111000000101101001010110110110110110011111110100010001010001100101110001011101011111100100010101111111101101011110001001111101111011100001111010101010001011111001111001000110101100001110001000010001011110111101110001110101010011101110100111110111010100001101010110001111011001101110101100100110110000000001110101011100001110110000100000010100111000110101011001110011110110010011010100111101001010111011011110001111110001000001101011100110001101001011010000000110110000101000100011001111011101100000010111101001101010111100000011011111001001000110100010010001011010000010001000010111101011100000001110100010000101000100010001000100101011010110111000111001010111101011100001111000000101100110000101010111011010001000111010101000100010011110101001100111010101100010001100101110111100011101100101100001000010010010100001110111100110001010101111011010101110111001011110101010101000000011011110110001110101011100110100101001111100011101000010011011000100001000100111011011111101010000100110100000110000101011101111100111111010000101110000001110001001001100010000011010011010111100110011010101010001100010100100110010110010011100011111001001000100100001100011111110110000100110111111111100000010100001011000011100100010111110001101100100101010101010110010000100001001011110100000001111000010100001010100101010101000100111111000100100000111010000110000010000101001111011001000001000010000101100010011011001110110111100001001100111011000011101110001000100010000010001110110110111010110000000111101001010010110110001011011100011101011101111100101110010001100111101001001011110011000110011110010101101110111011111100001111100010011011010100101000110001001000001111001010100111011001100110111101101001100001001000101110000001001111101010110000100101101010010110110001100000011111011001111110000010110010101001001010101000011010110111001010001100010001111010110001001000101011010100010000000101111001111100010011110110111101010110111011111101011001001010011100111000100100110011100100001111100010110001100011100001101011111110001101000000101111111000000011001000010011110001100100111001001011010010110111110010101111100101111001000001101000011001100111111100000000101000100001010010010110001110100011110001110000010010000111111001100001100000000111011101001111010110001110001111011111010100110000010111010101101000001011000111100010000010100111001101111011010011000100101100110100010001110010011011001101100011111000111101100001110110001000100101001010100000010000011100111011011000000010001010001100000110001010101000010001010000111000110110011110000110010000011111101111010100011011000001101010001111010111001001111001110111110011001011001101001111100000101000101111001011110111111100100101010111000000000111100010000000110011111000111010010110111001000010010000010100001110001011011111000000010100010000101011100100101110011100101011011100000100001110110101010010000011100001010110101000000011011111010010011000000101110101000011110110000100011100001100000111010111011000000101100000000100100010100100111101001011110101100100111101101110000000100111001101010100110100111110110100111001110000101000100001000111101110111001100001010001100000010101000011100001001001111101100010010100001000001011010101100101111100000100010011000000011101001111000001110101000001001100000111110100101100000001100010001111001100110101001101101010000101000011011110000101100111011110001010011110010001111110000001000000111110011001010001111001000110001010100110011000001000100000001010110010101100101111001101101010000110100101110011011100001010011101100000101001111011000010010010001110100010111110011010101011010001110100001100000001100011111111100101010110101111000010001000010101011111101111110101101011101100010000101000110111010100100110010111101110010001011110001101000110001110001100100001001010100100100011001110001011111100010101101111100111110011010011110111110010011010100001111101100000010000111001101110111011100000010101001101011110011110111100101111110101101011110010110111011011001001001010110111101011010001010011110010000011011101110110011110111110100101000100110100100010011100101000100100111111100110101100000011110011001100011100010110101110101101101000010111000011001111110101011110010100011010110000100001011101101000110100000000001001011010001010111100100000111111100100000010100111001101111001010110000011100111110101111010000001111011010111110101001001010111011101110000000100111111011010111101100000010010010010111100100000110001100010001100110100100010111110110111111101010011010101010101010011110000100100110111100110100010111110010010110010010110001000101011000101001000010111111110011100111011101101010001000011000010101010010001011111011101000001001101010010110001001000111010000110100000111110001100001011011100101101110100000000010111010001110111101011001101111100000011011001100000011000000001110001111101100000011001010101011000111101100011110110101111000110010011011101110000010111100010100001110101100100101010000001010000100000100101101101000110100010110110011010011010110110010011111010101000100001001110010010110101101001101101110000001000101001111000101011101001101001101101000011101011000101000101101111111111110100101001100100101111100001111011110000011100100001100000110011101000010111011110001000111100011000010110000100011101110000010010010010101110110011110010000111010110100101011110110001111000011100110010100100100010111011011110010101010001011000000110001101101101111101110001010110011111011001001011011101010011000101101100001111110000110000100010110101001011101011101100111111001100111001101011011110111010011001111010110111111111101111011111010010111110011111001000111000000010000010110011100100011111100110011001000101111001000100111000101100101001100010101101101111111111010101000110101010100100000001111101111001001000111110101010101110001000111011101001101001111001100000001010101100110100011010011100001111010011100111101100101101001111111010110001001010100000101110101100110010001101010100100010001001100011001001101111110001100101101110101011010111000111001000100100111111110000011111000010100101010001001000011011010101000101110111000000100100110100011001100101111100001100111101001100010100111111000101011000111001101011000011000001111000001010101111111011101111101010000000000100001100101101000111000010100010111111010110001101001110011010110111100100111001010111101111101011000111001011110110110110011010011110010100000001111100101000101000101001111101010101011000101111101010000011011011111110111010110110010010100101010101110101110011101000010111100100100100110100101111110110101110000010011111110010110000000010000101001111101111101001100001010010111111010011001000110111011101001001111111010010100101010011010101110100000100101111001100111110110111111010010010010100001110100110011111000001011000110011000000101011001101001011100111010101011000010110011010110110011101111010000111101011111111000010010011110111001101000110011001101101001111010000110000111010111110011110100100010100111011001101100000101110000100001101001110111011100111011001101011001101010100011100111101110111110010000011100110011010100110000001001000010101101010000111011001011010111001100100111011001010101000110100100101100100011001111011101101110110111001000001111111001111000110011101111001001110111011001110101100001011011100100100011000010001001000010011111011110010001001001000001010101001001011010011101101011100111010101110011000101010110101111001111000010011001011010101111111011111100110111010101001111110011000000111001011110001101111111101100100100110110001000111000001010100101011010011000011101011100000101111000111010100111111011011101100011010011101010001101001010100010011001001111010101011111110101101101011010100100001111010010101100011011100100100111101110000011010111000101111011000101101001101111110011101001001100010101100101101111010111000000100001111101110010000010100001100110000100001101110111100110110011010100101011000001101000101101101111111100011010111010101010100110100100110100011011100101000110100011000011111011111111000010111000100010001000011111111001001000110111001101010100100101110010101010100011001100001010111101001100001001111111111011000010100111011110100001110010100110111110100101110011010011001000001101100100010101010010100110101111000000100100100001111101101110011001101000010101010010111111101010010000101000001100111010110000010011111110110101010111000101010110100000110001111010111100000101111100000100011101101011010101101101110010011011011111111011100011001011100010011101110100100110011010000000010001100000001110110000111100101111010101001000100111001001101001011101111101011111111100101000011011100001101010011100101111110101100100111011001111111011101100100000001011100101000011110010100110111001011001001100011011100001101100001011011101101010011110011011001101011100110000000010100011100010010100111001101010100100110111111011110010000100100111001111010010110110110001111100001000110011001101100000101101010100010000000010101101101010011000010011101111010001111010001011011011101001100101100111001001111011011010110001010101000011001111101110011100110011111000000110111101110000100110010110001101111111011011111110100001011110010100110011010010110101001010110000001010011101001111000011001111011010010010010110001001010100010100101110010011110010011110011010111101010101100001101000010110010001001110011100011111000101111101010011000011010000101101111100011001011100001110101111101111001000000000100001111010110000110000111000110010111001000000111101010100111101010011101011011011110000000100000000010011000000000000111101101000011101111001001010011000010101100111111101100110100111100011101110110101011001100010010011000001111001110010101001010111011111101101000111011001010000011011001001010100001010000110011110111101001100010111010101101100111101001111000011001000100110101010101111110100011000010000110001010101000101001100001001100111110110111100101111010011101011000011110101010000011010111110000111001111001111001001101101000111000011111011100101100011001010011111100000110100011110010111110100011100111011011111000111010011000111010111011011010110010011100110101101100010010100100001110110000111111111000100011000010110011010110111100001110000010111110101010110000000110001001000010110001001111100110000100011101111100001101010101110010101101101110000001010111111000101000010100011011100011001011001111111110000010100001100010100111001100110110111001011010101001111011011000000001000111001011111111000000001101100000000010111010011100101101101100010001001010110111101010001111011100100000111110111011100100010100000111100100111011001001001000111101010010110010101100001000100000010111110101110010010000000001001001111100000110100001001100100001011010000010101110100011000111000110000011000010100111000111100111010100000010101110100000001111100011110101011000000111100110011001100010111100001111010000101101001110011001110000000111111011001000010101010111011001101010100101100110001101110101001111101111000110100000110010001001100110111110100000000000100110010000101111001010111000010001000000000001110101101110011100111011101100110001100100111110110000100111011111011111110111100000010100010011111111101010100011100110100010000010011110100110011010010100100011010101111110010100101011110011011001011101001100101111001001000010011111000001111111111101111010010000111101111010101111111011101101010001010011101000001100100101111100010000000111000111001111100100110001100111010010100000000111100101101111001101101110011101011011110110111101111111000110011110000100011000100100011011111010011111111010010101000011000110010001011111000100000110100100110100100110011011100111100110110111010001001110110001101010111010101111101011100010011010110001101100100110001101000101000110010010100100110000010001001111000100000100111000111101100010011010100110101111100101100100110011100111010111100110110110110110001111100011010001100101100010000100011010000110100000110111110011110100100111111011100010001100011100101000100001010110110011000001000100110001000000011101010010111111111101111111100111010101010011101100111001101111010110011101010011001010011001100010001000100010110011110111000100101010100110100100000101000100110111110001101010110100011000011110100000101000110111010010100100100111101100001101001010101110111110100000101011101100000110001111001000100101111011101110101010101011101011011100010101110100010110101110011001111011000110001011110011011010000011010111111110100110100101011000011110110010100001111111000110100000011010101000001010000011101001100111001101100000010000111101110100001001111000111100010001100000011011001101110110101101011011001010011000101100001110110110101100001001000101011110000110000101001110101000000011011111111101101101101111110010111000010111101010111001111110100001101110100001001010110110001001110010010001010110101100111111010000011000101011110101111101000000100110000111111011011101100010011100010110101000010011010010101001110001110011001010111110111101111011000100101000101110110101000111011110000011101010111101100001101010000010011001110000011110100011111100011000011000010000101101000111111001100101011011101000010001110111101110001010001100100010000001000101001011101000111001110010111010011100111101111010001000101111110011011000011101100001011011101110010100011100011011101101101011010000011111111111101000000010101100101110111010101000011111011110011010110010100001101100100100110001010011110101101101110100011011000110111100011111011011001110000110101100100001011100111001110110011101110101110010111001001001111000010101010011100101010001100000111000100101010010110111000111100010100011110000010110001011001100110100110100111101101101101000111001101111001101000000110110110011001101011010011101110101100100100110100111110001110100011101000001101011101111010110100100110000011110010000011111111111001110110110111000011001011111000000100110011110101001010000100010111010001000010111111111000110111111110101111100010110100010010011111000010110011101111001110000000010011000011111110011101101101111111000011010010011010000101110000111010100110011000111101011111111100011101101011110100011000010100110111010110001110000101011000100011010101110110101111111010101110000100000001001000100001110000111101100110001011100111010100111001110011000000011110000000000100110010010010001111011100010111011101100101000001110110100011011100100001001110010110101101001011011001101110101111110110110110011001000011001111110011011001001010100110110111001110101100110011001001101011100001010110000101011000100110011011111000000100101110011001111011001011101100111001111101000000000010101101111111000101000111010001101010011101011000100011101100111011100011011011011010011001011111001100010001101001100111111011111001110011101001111011111101010110100101100100100100010010000100110010010101000010101101011011001111000000001101100100010001011111011000000001111001001100010110111010010100110011110000001000010000000100001110000100011101111100111110010001001001101111000110010001010101100011010100000100000000101100101101001011111100101100110001101011110110010101101100101010010001101110100100110110001110100011001011001111010011001010010010001101001011010101111010000101010100001011111101110011111011110010000011110110001110110011110101000111110000101101000011010111101001111001100101010001100011000011101001000100011001101111000101011010000010000001010110000000110011010011001011101011000001000111111010010110111111011001001010110000110001101100000000100010010101100001100110011010011100111100001011010101011111110101101111111111110110011111100111110010011010101001101001010010101111011000111101010110100100010100011000100000000000011100101110001101000100001000101110010010000110110100110010101000001000110111011011011100111000101101001110100111100011001011001000011111101000101011110100000100010011001101100101110010000111010010110010101101111000100100001101010110111100000110011110100011001001000100010010100000111100010010010010011111110101111110010011001100011110011111101111000100101000011001100110001001001101110011101001011000111001101011001010110100010000010001101100000001100000111101100001100100101011011001010101011011101001101011000101110001010100011111010101011011001001111100110001000111011011101011101001101011000100001000010101010101010111100100000100011010011001101001001000010010101000010010000000100100100110001110001001100111110101000011011100011000001111101110101010011000100111101010010010010001100011111111101100001011110000000111110011100011101011110100111110010100011110110101001011010111000101010000001110110100111010001111100110111111101001111010111010011101101001000010111110001111001111000001000100011000110011010100111110001101100100100100110111001011110110100001111001111111100110011111001110111011001111101110001000111010000010100101011100111111100111110001100011011001010100101100101010100011101111110100111110001011101111111000011011010101010100010011100101011101100100011100011100010011001011011111111100100101101110111001010011100111000110111100111111100101000101111111011111011100111010111100100110000111001001010010110001010011000001110111110010111111011011001111011100111111001110100100010100111010011111101011101010001110010011100011110100010011000011100111110011101000001000011110111100000010010100111100100000111010010000101100000000000101111010001001101101110011000001101001010010001010111011100011010110111110010110001101100010001111111111001100010111110011011010011001000101101110011110010001010111100011000000100011010010001100001001101011111111101111100011101110010101011010010111010001100001000100001010010011010110110001100111011110010001001001000000000000100011000110000000011110001101000110010011011100000101110110100010000110001011110011010110110101110000000100001001110001111010011100011100100011111011000001010000010100011111101000010010010010001101110001100110000010000100001001110010110111110101000100110110100111011110100100101011010010111110101001010111000001101111010101011100010101101000010000010110111000001100100000110001101110110101010100000001110111001010100011101100101110001001111111011110101010000100000100001000101111101100111101011110010000001101101100111011110111001011111000100011010101010011001110010010101010110111111010000111001011100100001010111110001110000101011111000110111000111000110011100011010001010001001110100010111011001000011110110001101110000001100110110011100000010100010010011111110001110011100001110011100001100011101000100111100111110100110110000110001011000100001110111100001100111111000011000110100000101101100010111001111101011011011011110001010101010111011011000010111000010100101101011010111011011011000100110000001000110110100100110011010000001011100100001000101101101000100111110100010001111000010111101100000001111001001111111101001001111011101100001100111111101011100101111100100011100000111111001000010100001111111001011110000011000011110011110010111000111001100110000110010010000000000101001100110101101111110000001110011101100110011000001110011011000101001110010010111111001010110001011011111101100010101010100100001000001100010001111110011111111000010111100110101101010111101110011100001101010010010001111101011011101100101010100011111010011101111111100100101100010011011101011001010000010110101000111011000000100000101000011011010111101111010101101101100100100110100010010111110111100011001111011101101110010001000001100001010101100010111110110101001001110011111111010000101110110111011101100101001001101100101001100101011011011111001110110000010011011001111000101110111111000111010000110001101111101111011111011111111100110111110111011100000010011111011011000101001101010001001100001010110011100111000001110011111100101101011110101101011000101000010111111110000010110011010100000100010110100000101111000101101111010100000001011111101111111000111100011101001011000101110101010100101100110010100000111010111101011100001010111110010000011010100010101001111111011001110101010100001111011110110011110010110111100000100110110011111001001000110111011001010110111111101101100010001011100011000111010000001101111100000011000110111011100000110110001111010110000011001111111101111111001001011011011001010110001000011010110101010011101001001011100001110011101100101111110110010000011101100010011101110100000100110111010001110101000010000011010110101100101001111101000101110101101100101110101101011111100101011010100000111111110000100010110000001000101000101011001101110110111100100010101110000001100011001011111101111010010110101110111110101100010001110000111111010000010110000100000111101001111110001000010001010100110010000100011010100110110111000001110000111000100111100000010110110111000011000110011000100100011010000101001100001010101110001111001000110001010110110100000000011111010011000101001001110101100011000001010010001011110111000011111111110110001010011010011001000100101100010001001010110001101010001100101000100001000000101000101111101011101010000001111000110001011100011111010010010001101000100010011110001001100000001110101010101001010001111111101011110011110100100011010011010001111000001001100101010110110111100111010011001000100001111100001110011110010111101100001111010110101110011110101010101010101011110111111001111001110100110110010111100111101010010101010100011100110101000001010000000111010000001111000010101101101100100100101000100111111101101100010111101111000010000011101011000010101101011100101110100010011111010010001000100000001111110011111010110111011010101110101111010110011001101100010001001011100100111010010111110111101110001111010001101010101111110000010010011011010100110001110010110100111010101100000101110001101001101000011110001000110011011000000111011000101001001001010110111001001100100011010101101010010100111101100101110001100011100110001101011110111111100111111011101100000001001111100110010010101111000110010110111110111110011011100001111011100101000100100101001100101101001001001000110101101011100111111000110100011010101011001011001011100001000100101001110001000111011001111010111011100101001010111001101100011111110101110110011001000010101011111110100111010001010100111100000000001001010100101001001110100111000001101000001000101100101010111100010011110001110000110110010101111000100111011010000110100000010100110100101101110001100100111101011100110100000110010011010110101011100101000010101011010101001111011110110100001001110010110010110000000100100000001001011111100011000001101001001111010001000100111101010111100101111100110011111100011010100010000011000100111000010011000100101100111100000000110100111111000001000110111101101110010010010101011110011000101000011000100111111110001101000101100010101001001001101100010010011110101111011000111000110010101011100001100101010001010100011011101000001110100111000011001010101100011011011001110001011101001110010000111101010100010011110010101101011101101110110101111001111100000000010011101000101011111101111110011010000001001010011111100111101001000010111101010111011110001100011011011001111111000010110011100010001001100111101100010011111100110011101000000011111010110011000001111111101011011000001000001011011000001111000100000100001110101001100110010111010010011011100100011011010111010100110111100000001110110000011000110110000101001100101000100100000101110101111110111000011000110011000111011110001011011101011110110101000101111111011111001111100110011101110011001101000010110011100001111101100110001001000011011110010001110100101101111100001100000000011111010111001110000100001111101010010010111100101101101100110001010001010011001011001110100101011101011011001110011001000111001101111110011101010111000010001000100111010001101010010110111011111000110011111111001011000010100010010010001100110110101110101001101010001001111100011010001000001001000011001000111010000010111000001011100000100110101101000001010101101110001110001001110011011001000001101111100010110111101110100110110111011100010001011011001010011011000011111111001011011100010010011010110100011111100110010110011101100001001011101010010011100011011100111111011001000100101110111111011001001011111001100110110110011101101110000000000011001110111001111010101100010010001100100111000010110111101100110101100000101011110100000111111101000001101011001111010100010111000000111001000010100111011110101011000101010100010100111011010100011101001101110001111111010111011111011110110111011000100011111000101111010111001111111011111100000001010010100001101011100101101111110010100011011001011111010010001011101101001110101110101011100111001011010101111110010000101000001110001110010001111110000111010111110101100111100001000001111101011111000100000101110111011011001011010101101101111000001011000001000101001000100100001100000111001001010011000111001101001011111111100110111111001100001001001010010001010111011010101011011000111001010111000011110001011000001001111010110010100010011100100110100110010010110110111101101010101001001100010110110000111100111011000011111001011001101101111001110010010110010010110101001001100010110011100111110110011100000010000110111011110111101011100000100100101010100010101100101011000001010100001111101011110111001010101110011001111101000011100101000101100001010100001111010101010111100100111111100111000011101110110100110100101100010110101011010001001100010010001100000010001101010000011100010110110010000100010110111011101110011111111001101101000111001111000001111000011001011101100100001011001010010000010001010001000110011001111101110111100010001100111110010111111001110011100001000001000101011010001101001101111000001110000010011001001001011101000000101011110110000100000101001000001011011100101000000111111100011110100010101001010001100100001000101001100000111011001010010101011000101001101110001111000001011001111010111100011001000000001010000000001001001101101000111111111011011001101011101000100111101001101010000101110011000001110011010110110100111100111111000100001011000101010011001000110111000010001100011110010010001110100011000111010011000000101101001011110011110011111111100011000001101010011100110111100010101101100111001101101101000001001100111001001111111010101101110101110110101010110000011111010100100001010010000110000101000010110101100111001110111101111001010111000011101010010101111101101000100111000000001110110001100101000011110111011000111111010010100100001101110001010011010101001001101101010100011101110000010000001011001110101001110000110110100101010100111100111111010101111101000110000100010110110111110110101111100101100100101111101000001101000110101100111011011110000101101110101010010101010001010110000011101001111110011100010101011110010001011011011011100101000111101001001101110001100010011011011001101001000111110011101111100110101000011110101101100000100000011001110000100100001101001001011011000110101010111101101101100010100100000101000010110011010010101010010011100010010111110101000010100010010100010110101010011001101001110101000010001010110010001100110000010011010100010010011100000110010010101000101010111100010001001000010000010110011000011010011010001110111000101100001111101000100110000101110100001010110110010100100111011100101111110011111010100101011100100000101100011010100011111101011011011110001101101000011101001000111101100011101111011100111000110111100001110000000010100101001011111000101001001010111001110110111111111111010111100011111101100011010100111000110100111000000100100000100011101111001101111101001111010101100111011101011110000111011001100110101101011111010111010111110101000101010111011001100000100100100001010010100110100101111011000111111001000100011010110100000111010000001101011100010111110110011001100010010111011111000010110010100100011110110000110000101001011010110000110110001110111111110011010111010100100100011111111110010110101010011010011001100111000110001001111110111001100010111001101110110111101100101000101111000001101110000011111010111110100110100100011101011100100011001111000110100011000101110000010001000111100000000101101001110011110011110000010110000101011001110011000001111011011111011001111010000001010111101001000001011010110011011010001100100000111110111111101010000000100001111011110001101000001000010011011111011100100000011000010010010111001110110000110111010100011011100011100000100011110010010111100100100011001011100111101110111100000011010001111111010010001001111011011110110000111001101110001100101010000001110100000001010001011010111110001010001101111101110100111001100000010110110110110010101010101011010010110000100001010101011100111011110000011110101001100001100001100100100011111100011111111011101001010101011010000011000100110101011111001110011101011101010111110000110001000010001000110010101110110111000111011101011001001101000110000100000101101101110000011101101110001010000111110001000011010101101010101101001000111111011010011010101000110000001111111100001110001001101001011001100110001011101000110011110010011110010011101110101100100110010111100000001011100101110011000011011000010110110110010000111101001010001111111100010010111001000110000000001000111110011101010000001001101100111101000000011011101100010000111010110100011000101111011001011010100111011011111111111111010010011000001111010010000100010110110110000001110111010101001111110110111111010100110000000001100111000100001001000110100000101001001101111110011100011111001011001100011101111101101101001101001011011001000010100101110010100100000100100100001010111010111000010101111100011001111111010011100000101011011000001011000000011101101010011010110001001111100101000001011010111011001000000111000011010111100010011011110111101011011101010101110101111000110111000110111111100010001010000010011110001000000000111000001001000001001011100111010011101000110110101010110111111011011000111111110000111010001000110111011110100110011100111100111011110011001111011110011101101001101100011010100111111010010011100111001010111100001010000111000100010010001011000001110001001010111010001010010001110110000101101001000111100100001101001111000010110100111011101001000101010111111000111111001111101101100101110000110111000110110001111110010111001011110000000111011111111101010100110001001100010001000110110101010001011011101011010100010010111101001111001110111000000100101111101101110111110100111001001001001111100010011111010111100011010010100001101000100101000101101111100010010101011011111100100100110111110010110100110010001010010000111000101010111110101101111100001111011110001000000000011100101100111011101011000000011011000011110100001110001110001100100100011000101011100100010100011111111011000100010111110010100100000010110100000001111100001110000110000010110010010110000101101110110111001010001010110010111101000100110101000000010001001110001001000101110000101000111010011000000010101111010011010010000010010011010010111010110000111110101100111100100111011101000101011001010100111000000001000110111101110101110011101101101011010000100000000101101110101010010111001101110011010000111111001110011001111001001101011011101100010010100110101110010011101010101001011101100111000100101001001101110110111011110100110001100011101011111110000100110000100101101010101011111101000001110110110100111110101000001000011101100100000001101110111011010110001100110010100000001111100100101110011011110001101011011011101010100011111010101101101001011111001110111011111011111001000111001011110011001100110100110110111001000101111000111001010010100101100101001010100001001100101100010110100101111000001111001001001101011011100010101001010111011010000110110001010101111101011111111001011000110110000001010110101100110010110101010111000110001011110000010001010111100010101100111000010110111100011110111001001110111101101100100100011010100100110110111101011011001011111110001011101110101110011101110011101001011100101110111111110110110011100001101010100111110011010110010010010101110110101100011100001100001001111110100100000011111011100111111011111010000001101110000100101010110010011000110100101000010100100011110011000110110100101100100001100000011110010100100010001010000000110010010010111101111010110111110101001001000001000011111001001101101111010110100000001000100101101100111110110011111000011111111110110000100110000000111010111011011101101100010101100011010101001101011111000111111001011011111011001010010100100011110001011100000001011100010110011010111101101111111111000100100100111100111001110100111111101101000010110110111111101111110001000001000110100000100001001011000011000110000010010000010001011101110111110101011001101010111010110011000100101001000000011010101100000110100010001000001101001001111110101000101001110000111101110010101001011010001111101101100000001100101000001110111011111111000101101101110110110111110011010010101100010001000100100100000010001011011000101010100000011100111000100110100011000111010010100101111111110100000011101101001001100100101001010011010000001001010110010011011101101010010010111000000011101110110011010101000110001011111100101010110011011111101111011010100011101000101000010001011110011111000101001101110011001000001111011100000011101111001011101011001110101100110011001001001101100110110000010111101001010111100111101001010111000001010111010101110100011010111000001111100110101100110101100100011111000111000010110111110011101001011011110110011110110110000010100010101100001101111100111111111011000001010101111110111001000011010011010110111100000000010010011100010010000101100110110100001000010111011100010101000100100001011110011111110000010001111101000011010111001010101010111001011101010000101110001101111010011100100111100100000100000001000101011111110010101001100001000000011011010110110000101011001001100011010010101010101010000000110011011010011011110011011100110010000111010100101110101110101100100101011100010100010101001000011010100111100110111000010111010000101011011000011011001100111000100111111001100101101101110011010110011101011101001111001111101001010010010011110110100110101011011010011000110001110110100001000011010011101001011011000110100011000111110000100101101010011000100000111100101000101010101001000011011111010001000110001100010001101010110100010001110110011101000010010110001101100000001001110011100101000011101000011100010001111100000010100000101110010000000001110001111110000011011100101101001000110100001011000111001110001011010010101111000111000100101000100111000110001001011001101011100111100101100010001010011110000100000000011011001001111101011100101001011010111111000001111001100001110100011110011000010101101001101001010010101000001101100001000110010100110110100010100011110010111001010100100010010111010011000010011011100100110110011111000011010111110010001010101000111100111010100011000001100010110111001011111001010110100001011110110100010000111111101101000011100100111010110001000001101010111100011111101001010110110010110101010000010000111010101011110101000001111101010100010100100100110111101001100111000100100100111100110001111111010000011001110001010001111010011111100010111110011001110001111100111000100011110001100111111011100111010001010010001110000010000100010000100111101111000000111011000110001111101001111101111111111111000110110111001111111011100011101001111111110001101000001001101100110011011111101001111001110000101011000111100101110110100000111111000111000011111101110000101100100101110010001001011110101111100101001100111101010110111000001111001101000011100011110110101100010100001010100001101011011111000011100100001000111010000110011111011011011110100000011100010011010100001010100111100110111100001100110101110110110111001010100110000001000000000011011011110111100000010100111101011010011001010001110011111100101000100001101110100011010100111010001110010000000000010111011000001111111111111100010101111001101010010110111011100001001010101101011100110011111001101010111010000001101101111000110101001000000100001111001100000000000011111111110110111111010010111010010000100111011110110000011100010010010110101101100100100001001110011111101111000000111010111101000111011100100001101001001011001010111111001001100000000010010100100100010011011101011000100011111110111100110001011001111000100001000001111000001100111010001100010000000101011110101111000100000101010000000101011100110100110100100000110100101010010101111111001010011100000001101000111010101111100010011101110011111001101000000100010100100111100011111010001010110100011000101100100100100001101000010110111100110100010010010001010001100011101111000001011001000011001100010010111100110011110000001010100000001111000101010100101101100011010001010011011000110001010000100010011011101100010001101100100000001000110110000100000110010111001011010101011000101010110110001010010011001011101001001101101000111101011001011011010001111010000000111010111010101110100001010101000010100001100010000000010010000100000111010010110100101111001101001100011011000100000111101000010100110011101100011101101100000111010111000000111111110100110111010100100101111111110001000011101000101111100001111101000110010011001000010001000000001000101101001010010011100100110011010001010010010111011100000011100101001100100010010111010101001000101001100010011100000010001011100111000100000111101000010000101010111111101111001001100010110101011000010110011100110101101110011011100010000011001100001111010011101111111010010100101111111100001110011011011111000000011011101011010001011111001011010110100011001101000101110111000111011001000010111000101001101001111111111001111101110001001111010100101001010001010011110010011101110111110001101011001001001101111000110010001101111001001111110110000100000100000111101011010100110010110011100001100110100101111001111001001111110000011011101011010001010010001010001100001011000101110101001110110000101110011010010000110010100010010001011010001100010001010011101001000000010101100010100010110010101000011011011010110101001011001010111111001011101010010100101111110000000100000010111111100011101000110011000011001001100011010111010010111100111000000011111111101111101001110010110111010101101001111011100111000001011111001010100000001101100011010101000100011000110100011011001011100101100001110011000011101000011000110001010010100001101000001001001101001001111011111001100011101111010110110001010000001011111010000100010000000101000001010011001111010010110111010011001000000101110110001110101101010000110110001100100101011000101110100110110100110001111100011000100110011000011100100000100101110000010100110111111011001100101011100101110000000010011010101101101101010110001001010101000001100001011110100011110100000000001100010010001110111111010111010101001100001010011111011000000011110101010100110000100001110010110001011011001011101110110110100100100111001100111011000001000000100011001101101111000010000011010010001010011010101000011011110011110111011111010110101101101100100101101101100100100100001110101000110110100110011101010010111110111110011001110111111101100001010011101011010010110011010001101011011101111010100110000010100011001001011101101111100101111011011110111111100110110101111000001011010011110100011000101001101100011100101110001000000000010001010010101011001011011101100010111011101100001011100010010101000011101111001011111111110010100111010001111000000110001101101000000100001011000001010111110101011011000100001000111011101011111010110001001010010011101111111110111101101110000111111011010101110011110011111110001001000110101000010101011000101000101111111100010110001110000100011100010100011111000000111100111110011001110010111110110110001011000001110100100011000000010110100101101111001001000001001011001010111000000110110001111010111010100001111100110001010001101101110011011001111011000101010100110100010110001001111011110100101111111110000001111000111111100011110101111000010110111100000011111101010111001010100101100101110100101010110000110010100110110001001010001100110111110110100100001011011111100010111011001011011011100111111111011001110001111010000000010101110010110100101101011001010010010100011010010101100110011100001101100101110000000001101001100101011001111011100110101100100000000101001011101001000110101000010111110110000111101111111000111110011110011011000100011011101011101111001010101110111010111110101011010011010110110000011000010011111001010111001100100100110000000011110001010100011010010111100000001111001011110010001000010100111011010110010000001110011000011000100010111010010001000010100011011001010001010101100100101001111011000111110000000110111101001101101110000110000010011110011111100101001111011101100111000000000110011110010000100010001110001000001100001100010011111111000110110111110110101111001110100111110011000000100000011111100100101011101110100110001000010000010100000110000100010100011110101011110111111100010011100000111000011101010101110110100110010100110011101001001101001011011000111100011110101000100100010110100000010001111001010011011010000011001001011001111010010100011111101101010110110100100011101101101111101010010100001110100111111111000110111100001100100011011001001101000111000011110010101011011110000110111110000000110010001111100111101101010111110010001001010110110101011010110111101010011101001110101110001101100101010101100011011110001010100111101010001010110011101101010110110010001001110011111101100100110010010110010001100110101100110101010010010001001100110100111110111110110111001111111100101100001000001001110000101100010001100111001101111010000000101001010110111000010100111111100000001001011101110110001010010001000011101101010010011001001000101000111001110101111011111011001100101010111000000001011111110011010011001111011111000010011001011001011010110010101001010100101011011000111100000000011101110000001100110000011100100110100101100010111010011000011111111100000000010110111100110100011001000111100111111010111110011011101000010011111110100101011001101110011000110110011001100011011100001011000111010110111010011101111101111010001110101101111101001000001111011100001111000001101000101100110100000000001011110010111011011101011011111111010000100000011110111010100000111111000010110110111110101011011100101011101001010011010001100110111000111011001010000111000110110001000101001110111100000011000110101111001100011001000111111111110111100001010111111000111000001110010101011011100100100011000111001110010010111110000110101111011100011011111110110110011010111001001101111010100100101111010001000110101100000000111001110001010100011010101001000000100111111101000101110101011011111000111011100010011011111010101000000100001001010001011101011000101000101100101110000001101000010100101111011101001100010111001011010101101100010000111111110010001110110011110101000000101001101100011111101101101000000101110110001101111101101110001100010010000100011111100110100111001101110001110101100110010100101100110000111111101110101101001001001001110101010010101000100111011011011001101000110011110000001001011101011000000111110111100010100101000111011000010101110010111110000111011001111001101110010100001101000111011110011000110101000111000010000100011100000000111110101001001100000000000100010110101100000111100011110101110010000000101111010011011010110011011100101000111010011010111100101011111101100010011111111001100100011101011110101000110001100111111010001111111111100101011111011111101001011010000110000111000100000110101011101000001111101101010001101010000010110100100010011000001100101011010000011000100011001110000101101010010101110010011010101000101100000000111000010001011011001011010110101010111001010110111001111100010110101110011011010110101010011011010110001101001101000011100110000010100101000011110011010111011010011011111110000001011000100010000111101101011111101001010101001001001011011100111111000010110001000100100100110110001110010110011110111011111001000101110101100011100101000101000001011100111010101111111111111001001010011111011111111111110001111101110110010001010010100111111100001001011010100110011000100110001101101001001011010110100000111010000111101001111001010100000110100111101100100110111010001000110000110000101000100111101100100100101110110011010101101110111110000000101110000110000001010010101010001110001010111101111001110101100000110110110001010100011001101001001010110111000111100101111101110100101010100110110001010111001101111001001011011110110101001100100000000111001111110011101000111100011000100110011100001100101100101010001011011110000010000100000001100000101110111100011001111110111100101010100011001101011110011111001010111100101000111101111000110110001011010101111101110000010111101000101100101011110101000110111100110011101010001100110000100011010010100000111010000010101110111011011001010010110001100101110010110101000101011110101100110111011111111110110010010111001100010001110100111100110111100111101000101110100011000001011001101100100111110010110111110110111011000000010010010101010110010100001011111011010011000010101110011110111110001110000110111010111100110101001001010001011010011010000000100001111101010110010011111011111010011000001111001011000011001111001000001001101100010101111001110100111101100010101000010010100110100000001101010111110110110111001110001010101110110100100011011100101010000001011111011100001001111000010011010011001001110001101011101111011001011100010101100100111010100001010001001010010101010101100110001100101000101001111000101011000001000001101110110110011101111001000100101101110000010111111011010100110011001101100111111111101101110011010000001000110100010000100011100000101001001001100000001000100000110111000011011010101111110011010001010110111011000010101110111011010110001101011001011011101001011101110010110010001011110001011000101011011100101111011100010000001101110111011010110000010011001110101111111110011001001011010001111110100011010000000111010111001001111011010010001010010101100100111100001010111110110100011101100101010010111011110001011111001101111010001010100100001000110101000001000100001010001100001100111100001101111101011000100001000010101101110110101111111111100011110011011111010011100010110010000110001001111011101100001101101100010101000011010100110111110011000011110111100000111101101011000001000010000100110101100101000111101101011111110110111010100110011100011111100101111010101011110001010100110111111010010110101000100100010100000010101100001101101101111101111010100101001011001101111010100111010011011101001101111101000011100100010100101110010110001100011001000110100111001011010100101110110000011010011010110100100110111100000100011001011110011010110010110101001010100001001111110100010101110011111011100001101110011001110001111101110110110001000100111111011100011001111011010100011101101010000110101010000001011000011011110100000111101001001000000111100001101100000011101110111100000000100110000001111101111111101010010100100001110101100111100010010101101001101001011011010110010010100100001000110001110011011001001010000110001011011000011001000000111010101110000110001101010111111001011001000001010100110000011100011001110111010011011011001100000111010011111010011011010100100110000000011010011101010000001111011011010001001110110111001100110100010110010111010100110010101001100101001000100011101101001100110100110001000111111000110010010000110001011011001100001101000110010111101101100110010011110101010110001000100011010011011101111101111110011001000111101111110110011111010010001010111110011101100011000011001110011100011110111011000011101001010000010010110100001001110001011100111101110111100000111110100101000111011011101000001011010101010100011111101000001011110001111111001010100111100011110100111011100010011000110001110011011101110000110100001000111111000001001001101011010000101101001110010111100000111010111011111000100110011001010101000000110110100110001110101010010000111110101111000000010001010001001000010011111110011011100011111010110110011011110000111001000111101101000110011000011111010011111000000101101011011010000010101101001110001001101000010111101001111010001101110010000100111101100011010100111011001111000101000000100110011000110100011110100000111100110111011110001110101100011001101100000101001101011100011101011010111000111011110100110010001000111001111011011011101111010100111011110001110100101101000011101010100101000110000001100010110110011100000000010011111110010101001110110000111100000111110000010001010010111010110100000001111000111011010110001001001001011000111011011011010100111100101001111001010101000101111110100011111001011000011101110101101000101110110110110110000111101010001101111000110000010000111110011011011001110111111100000001100111101101011000110011101001010110110000010101010101011000011010100100011010000011001011100011110110000011101010100001000101001111010010010111001111010011100000110011010110110111101101010010000000111111001110100111111001111110110100001001100111110000100101010111000001111001010011001010010101000010101110000101111000111111101001001011011101111111101010010011011000011010101011011011000110010011111101000011100101111100000001100000010010010110011011100001110110100010101001000100011011010000110100011011101101111010010100011011010000111000011101100111001000110000111011000111100100000101100000100100011111000001110011100001000000000001001110110101000010001001110100100110001010101000001001010110011001000100001100110100011011001110001110111101100010100100001000111100000101000010110011001001101100011000011110110001100110100110110101110010110110111110010110101100010111100001011101100011110011000100000111001101011010110111011001011100000000100011111010100010100000011001000100101000111100011000010010111010100011111010000111010001000010000100010000001111011001001001001000001111001100000011100001110111010111110001111000100110100010101001100100010110101111111111100000010000010001001100100111110110101110001000011101001111010101110110101101100010001111010101101010101011100101100000011010111000010110101010001011010111111101101000101011001110010110110010010101001100010110100011100011101111100011100000011000000010011000011011011101101010110010111100010000110001001011101111101010010111100111011111100110001111101100111011111000111011101100110001001000001000010010011100101100110100001011101000011110001010111101000101100011111100100101111011111000111110110010000010100001100100011000101101100001111100001001010000010011101110011110011111001101010000001000001000011001101010100101110100000011011011110110101011110000110101001010010001010011011111111010000101111011110001111101100110010001101101011100110101100010101001111101111100101111101001101101101111010000000010010010001011111110001001010100111100011101011100001000110101110110000010111110010101010111110111000000010100000001010100001000111100101000101000101110110010000100011111001101101111101000000011001100001101010101001110111000110101010111111001101001011000101100100101100010011010011011011100110101011011111110101111111000111011111000000001101110000100000001011101000101001010100111100110010110101110000100011100010101100001000001011010011110001110011010110110000111001110010010010100011111101001011011100001111101001011000010101001010100010010000111111100011011100010111100000000111011110101100100111001101111001000011111000011011111010010011010111101111101100000100111101111001110011000011101001011111111110000010110011010100101101011111001111010110110111111100000100100001110100110001001000011010010101111110101010011110000000001011111100000010010011000001110101010011100001010100000111101100110001111100011000101001111101011011000101001001010010000111001011001110000001011101000100000100111010011100111100011100111100010101111100110101100100011001000011111111100101101010111000111110110100000000000100111000111001011101111100110000010111001100100110110000101010001111001110001100011000001100111010000011100001110000101101010110111100101100011011010000000111100110110111100100101010001100000001001101010001101000100010111101011001100110111001001000110110100010000001011001001010001110000110000100000101000100001100110011111011010111010010010011110000100111001110110010000101000101100100100111001111010001101100110101010001001110000001000100111101001110110011010101111110010011100100101111110010010101100011000010001010011100110111110000010011110100011000110101001000001100001111100101111001001101010001101000100110001000101000111011011010111100111001011001101111111001110000110101111010001110000100001110001101011100101001010100110100100010011000100000010101001001111001011110101010110101001100011011101101100001001001000011001111101001001001110101011111000110000000111001110000101101010110111000100110111100000001101100100001101000111111000001010001111000010111011010110101011110101000111110110110011111101001010000001110011110100000111111001010001110010001010110111010111010010011111011110110000000001010000011011101111000010010101110100000000110100000110110100000110111011000011100001011101101011011101111000000000000011110011110010101011110011100010000111011110010111010101110111011000101000001100100000111011010101010011110101010100101000110010001101010110111010011111101111100101111101011101010111110010010010001101110010000100011110100010110001001101001000010010111000110100001100001100011000110101110010000000011011101100110101100101011011010111101011111011100010100001000001010100011110100001001011110111011000011101111000010100111011100100000000000001000011110001110011100000100011100111111110111110100010001000011100110000010110001110111010000010110010010000111100011111101010001000101010111001000010010111000000111111110010110010010001010011001010111000011101111101111100111001011000001111011001011011001100001110010001011000000100010001010010111001010001001011101011011001000000001111010011011110011000111100110110010011011111001000110100111110000100000011000001000011100111011001010101010100000010110011110000000010011101110101011111110110000100101101110001000011001000000011001001101111000100010110100111101001001111110011011100110000110010101110011011010001100000110111011101011011001001100111101000011010011100100111010110100111111110000110011110011110000111101010000000011010110011111101011010101011100111110110000000000010110010001100100110000001010001100100010100010010110010010101000100100110010011111001101000101111011111000100101000000010100000111111110110011100011010101011100100010100011011011011010111001001010110010000000011000011110011101110011111110100101111010100001110000111100110011110001110011111000111101000000100101101011110011000000011100100001000111100101101001100101101110000111100011001001010011010100110011011010011011101100111010011011111001111011000111101011010110111011101100111101110111101010110100011101100000010100010101110001000010111101111011111010111100101010100000010101000110001011010101111000001000010011001101000010011000011010011010111110010111101010011001000001000110100001001000011011000001100000101100011101000000001000001011000100110101010110001001100100110110111111001011110010111101101111001111101101001101111111000011100011010101001111011111100011111110001100100110101100000000001010011110010010101111001101110111100010101101111111010000011001010111100001110000011010011011110010101000101000110111110000001010101100111100010111111000111110001000111111011100011000010001100011001010100001111100000000010100110011110110111000011001110101001100000111000010011100010010101101110000101000110101111000010101101100001101001101110110101011010111101010111010000111111101001101101001011100110010101110101010101010011100100011100101111111101001010110000110110001000011000110111011000010000011111100010111101111111111010110100001000101001001011011101110110011011001100001100100101011000001111101111010010110010011000111101101010100100001110100000100111000011011010101111001001100111111000010110110011001001011010010011000101010101110101011101010011011101111010101100011010101000001011101110001011010100101011000111100011000011000011000111010111001011101111101000101010101011101100100011111110101100111000111010101100100111100100000111011101010111111011111001000100110011011110110011011001011100011011001101110111111100011011111000010010011010110100100101101011100111101011001101101011110101101101101100111101110001110010001101101010111110101010101101110011111001011111001000110001001001000111100111000111011101001000101101010101001101010001101010111101001011011110101101110011010010001100001001100010010100111011010101010001001110001110011000101100010001101101100101101111011011011100011100110010000011110101111010101000011010001011101000010111110010010000101011101000101011000000101100101011100101110111101001011000101010110111111010001111101010000110110110101011101010010010010010110010100001001001100000100011101011110001001011001001101110000001110001111110101011111000000100101001100011100011011001001001001111101010000000001110111100101000111110000100010001110000000100101111010010000100101101101000011101111100010100100011011101011010010101100111111010000000110011111110011010001000110111001101101001010000101111001101010110110000100110001101111111100011000011010101001011100011110001000101100010111101000100111000000111000001011011000101011000001100011000010101111001000100111101011111001111111001001101001010010001101010001111010110011101001010111011100101001111011000000001100101011010100011011100101000110010001111001010101111011100110010110101011001111100011100000110011011111010101010101010010001100110000111101011000011110110000110110110111111000111010101110011101100011001101001001011000001010011010101111101001010100010110110011011000101001111001101100011001100101001111011000001100100000011110000000111000111000001000110111000010100100101100110110110100001110010010110011010100000010101100100100100011101011011000000001001110000001010010001010111100110000101101111101010000100101010111100111101011110011100101111000111110110010111010110111010001110010100000100001000111110101001100001101001110110111101000001100111000011000100011100010101011000001000011010111100100100010011101000001011000100110111000101100000001010000000001101010101011110001101111100001011010001011110010010000101001110001101000010110110000101011111110100111000001100100010111001000010110101011001001101111100111011011101010011101111011101010111011100101110001111111000111001000110000100011100111011111101011100010011111011001000110111001011000000101011100100001110111110111100111111100101110000101011001000101110000100101000110101100011101011100110010010001101101110101010011011010001110000100010101110100110010101001100111001011001010110101000100111111110110101000111000011001010000001101001110001100111000101011001101010110010111100011100010100101001100100011001111001110010101101110101000110100101110011111111110110111011110110011110001100001100101101011101111101101101000011011101001011100001110011111101001111111101001110110010001000100010010010110000011111001100011011011110101111111110010111101101101111000010111011100010100001100011010100110010111000000111001010101100001000110111001100110100010110111101101110100000111100000000001111110101111010011001010110111011010010010010100011010010101101001001101101111111111001101101110100011010111001000110000010111000101110010010000011100011000100010110011000111111100100101101000000110010111101110001111101010110110010101100111101110011001011110000101110111100000101000101010000000111100000101001111010001100111001110111011000011110000100001001010111100001000100001101110000100011111001001011111001011110011011010111110101000110100010001110000001100101110101001100001110000011011011100101111000000100100011110000001100111110010111100010101100100000010000101011101100111101001101100000101000000000110111100011111101000000111011010011000000111111010000011001101000000110010010000000100111101100111111000011001111100101101000110001001010110000000011001010100010100010011100011011110110001000000000001011001000010000000111111100110011001100111110011011101000110010001110011111111100011010011010011001110000010110011001101100000110101011111000110101110110100100100011100011011100011111111101001000011011100101100111100100011001100000001110001011001001001110111111001100100000010000001000110101101101001100010111010000001011000000010101000010110101100001011001111111011101000110100110001100001100100011110101010100001101110110101110110110010001010001101101101101111010110111001100000101101001011111001001111100011010110000010001110100100000110011110101100110111110000111110111110011001110111111111101110011111010101001100110001000110101001110101101000110100100101001011101001001110100000010000101000101010100011000001001010111011011010101010111110101110110100101010011110110001101010111000000110000110100011101100101111011011111010100010001001010000001011001101101111101010000100000111110011100101010010010101000110010001101010110100111111100001000010011100100011111111101101110100001010111001000100101001110001000011001111101100111011010100100000101100101101110110100111100010100011011001000101011111110001000011101111100111100001011010001010100001000000101101110101100110101101100010000110000111111111001100011100011010010110101110000111111111110101111010010000100100100000010100101001100110010100101011000000000110110100011101111011001100001001001000000011010101000110000001101100101111010001110001101011101111110111110110011110001110101110100111111010000110100000110011110100000010100001001010110000001100110010010011100101100011101001000011100110000010011111100011000011001110100110111100111001001000110100111111111110101100110100111111000001110100001011101101100000010010011010110111011100001111010100010010011110001011011011010101111011110110001101110111110100010110001011111000000110011111011000101000010110010011111111001111101101100110000010110110100110110110111011100101001011000001000000010110100011000001011101110000000100101001110110000110111010110111011101110011111011110110110010010101101010000000110010100011111001110111100001101011001111110010111000111101101000110010110110110100100011010011100111100111101000111100000010001111011101011010000011001111011101010000011000101111011000111110101100101010110001100011011000010110010111010000000110000001111111100111000010010010100010010011101101101101101111111101011101100000011011101011111001100011111011111100010100000000010110011001000011111100101011000011000110100111111100010101111100000101001001011100110111001100110000100111110010110001101110000000011010100110011010001101110010100111101111000110110100111011111101001000001010101111001000001110110100011101011010111111011101100001001111110101000111101011001000111001111100100100110001100011111010111010110011110011000011101010110111110001000100110011000011000010100100110110110101101110110000111111010011110101111110010010010110001000000101101100111111001000101110101001101000101000101011111111101011100110111010110101111000011110110101110111100011110100011111010001010101111100000011010010010111110111100110101110111000010101010110011001110011001100011101110000001101111110000010011101111101011111000111010111010011000100101110111010111001110110011101111110010111000110100111110000000110111011100100110110101000011100011010011000000011111111101111001010000011001110000110110101110111101010011010101001010011110111000100001101111010111110101111100111000001110001101001010001110001001001111110110110011011101111001010010101100101011100000000111010010101001000010101110011001111100111011000011110111110111000111010011001011111101101101101000101111101100000000001010010101111110001110100000111000101111001011101001111011001000110111000100001111010001100101101010111011011101001101101101110010100001010100000011110100001000101011110011010000100110000100110010001001111111101110101010100101011110100101010010111010100000101100100011100011111010011010001110100101110010001110100111000101100000011011000000011001100010110011011010101111100100000100010000101011101111011111001010001001110001011110101100000000011110111010110101000001001110100011001000100110111111110010000010010011000110100110011111101011110110111001110101011010101111001111100011100000100110001010011010010110010110011101010000011111000000101010100101000010000111110000110000010111010010101010110100111101001110011100001010110000110101110100100001111101110110001011001101011011111110011111101101110001111100110101011100101011011011010110111001000111100001000100111100101100110101010111000101101010010011101111111000000011110001010010011001110101100000000011010011011101110011101010110101011111010101001010000000000110001101111100011010011001010010000101011110010000110000010101001001111000001";

	TYPE registers IS ARRAY (0 TO N_EVENTS - 1, 0 TO 3) OF INTEGER;
	SIGNAL registers_check : registers := (
		(0,0,0,35),(0,225,0,35),(43,225,0,35),(163,225,0,35),(163,225,0,23),(163,146,0,23),(141,146,0,23),(52,146,0,23),(52,186,0,23),(52,186,0,114),(52,186,119,114),(52,179,119,114),(52,87,119,114),(52,122,119,114),(104,122,119,114),(104,122,122,114),(104,122,122,186),(111,122,122,186),(0,118,0,0),(0,0,249,0),(0,243,249,0),(0,243,249,25),(0,170,249,25),(0,170,44,25),(0,170,92,25),(0,157,92,25),(0,157,219,25),(0,157,164,25),(0,157,247,25),(0,157,247,96),(0,157,178,96),(0,200,178,96),(0,200,240,96),(0,251,240,96),(0,0,39,0),(0,5,39,0),(0,5,39,200),(87,0,0,0),(87,0,1,0),(87,0,191,0),(183,0,0,0),(132,0,0,0),(132,32,0,0),(132,168,0,0),(132,168,0,141),(132,222,0,141),(132,142,0,141),(132,255,0,141),(132,63,0,141),(179,63,0,141),(100,63,0,141),(100,63,0,1),(232,63,0,1),(0,0,141,0),(0,0,141,59),(53,0,141,59),(53,0,141,130),(53,207,141,130),(53,83,141,130),(53,83,22,130),(53,83,22,21),(53,53,22,21),(53,38,22,21),(177,38,22,21),(177,38,22,219),(224,38,22,219),(64,38,22,219),(64,38,22,182),(64,38,26,182),(64,38,26,180),(64,87,26,180),(225,87,26,180),(225,87,26,113),(225,14,26,113),(149,14,26,113),(149,14,232,113),(61,14,232,113),(61,14,105,113),(61,166,105,113),(61,166,105,46),(61,166,209,46),(61,23,209,46),(61,23,209,76),(61,23,209,205),(61,14,209,205),(61,14,209,108),(0,0,175,0),(0,0,175,255),(0,0,251,255),(0,224,251,255),(182,224,251,255),(0,0,0,196),(168,0,0,196),(168,0,103,196),(168,0,103,167),(168,0,75,167),(168,48,75,167),(168,48,57,167),(168,48,57,221),(6,48,57,221),(0,0,194,0),(0,0,194,186),(47,0,194,186),(47,0,194,115),(47,44,194,115),(47,44,155,115),(234,44,155,115),(245,44,155,115),(245,44,3,115),(245,44,3,135),(245,44,3,19),(1,44,3,19),(65,44,3,19),(136,0,0,0),(136,196,0,0),(136,196,0,14),(0,0,0,213),(0,0,225,213),(0,0,225,8),(0,0,225,237),(0,0,181,237),(0,0,181,219),(0,0,9,219),(0,0,236,219),(0,162,236,219),(0,220,236,219),(0,220,71,219),(0,220,54,219),(0,0,54,219),(122,0,0,0),(184,0,0,0),(184,0,48,0),(126,0,0,0),(126,15,0,0),(126,15,0,229),(126,35,0,229),(23,35,0,229),(23,230,0,229),(23,230,0,76),(23,230,71,76),(23,230,71,191),(23,230,71,160),(23,230,123,160),(98,230,123,160),(98,230,123,0),(98,230,139,0),(98,230,139,210),(98,5,139,210),(98,5,139,202),(98,5,122,202),(98,5,79,202),(0,0,0,50),(183,0,0,50),(183,0,0,44),(138,0,0,44),(138,0,0,132),(138,142,0,132),(0,0,0,142),(0,0,3,142),(160,0,3,142),(160,0,195,142),(160,0,114,142),(160,26,114,142),(94,26,114,142),(94,26,114,236),(94,26,114,204),(94,26,114,139),(94,80,114,139),(17,80,114,139),(111,80,114,139),(0,80,114,139),(0,0,195,0),(0,119,195,0),(0,119,195,243),(64,119,195,243),(64,248,195,243),(20,248,195,243),(20,248,184,243),(20,248,209,243),(20,248,102,243),(20,248,238,243),(20,248,199,243),(20,248,7,243),(249,248,7,243),(249,120,7,243),(20,120,7,243),(0,0,70,0),(0,30,70,0),(0,30,70,3),(0,30,70,72),(0,0,0,47),(116,0,0,47),(116,0,50,47),(29,0,50,47),(101,0,0,0),(101,0,0,36),(0,0,0,38),(0,0,0,203),(0,0,204,203),(0,0,204,84),(0,30,204,84),(105,30,204,84),(105,30,207,84),(105,30,207,150),(43,30,207,150),(43,30,207,110),(43,30,96,110),(43,241,96,110),(43,241,40,110),(43,241,40,251),(43,241,40,38),(43,219,40,38),(43,219,41,38),(43,219,212,38),(43,170,212,38),(43,237,212,38),(43,36,212,38),(43,36,74,38),(0,0,0,185),(0,88,0,185),(0,88,0,231),(0,88,63,231),(230,88,63,231),(230,182,63,231),(197,182,63,231),(197,182,217,231),(197,182,217,160),(197,182,119,160),(197,59,119,160),(157,59,119,160),(157,154,119,160),(157,154,119,94),(157,154,80,94),(157,154,80,170),(157,154,80,236),(157,154,13,236),(157,154,23,236),(157,154,23,54),(212,154,23,54),(212,154,193,54),(212,87,193,54),(212,87,193,0),(239,87,193,0),(239,87,193,186),(0,158,0,0),(0,158,0,197),(161,158,0,197),(161,182,0,197),(161,182,0,93),(161,182,138,93),(161,182,179,93),(161,182,245,93),(161,182,245,98),(161,182,245,187),(161,182,84,187),(161,183,84,187),(19,183,84,187),(66,183,84,187),(66,183,216,187),(66,183,216,98),(79,183,216,98),(79,183,192,98),(0,191,0,0),(0,191,0,68),(57,0,0,0),(57,0,0,247),(214,0,0,247),(214,0,0,62),(214,124,0,62),(34,124,0,62),(34,124,0,128),(34,124,0,247),(34,124,18,247),(223,124,18,247),(223,124,33,247),(223,237,33,247),(223,237,182,247),(223,237,62,247),(223,237,82,247),(223,237,82,73),(25,237,82,73),(25,237,119,73),(52,237,119,73),(0,0,70,0),(0,0,70,179),(0,0,23,179),(0,0,116,179),(0,25,116,179),(0,0,0,65),(0,0,166,65),(0,0,166,34),(0,0,196,34),(0,0,196,91),(0,0,50,91),(0,0,16,91),(0,0,141,91),(0,0,141,239),(67,0,141,239),(67,0,141,17),(67,142,141,17),(67,142,152,17),(67,142,125,17),(246,142,125,17),(246,32,125,17),(246,32,125,213),(246,32,125,255),(166,32,125,255),(166,32,251,255),(166,248,251,255),(166,248,251,228),(166,248,165,228),(0,199,0,0),(34,199,0,0),(34,199,247,0),(127,199,247,0),(138,0,0,0),(138,9,0,0),(69,9,0,0),(69,9,86,0),(69,1,86,0),(69,66,86,0),(76,66,86,0),(76,66,86,168),(100,66,86,168),(100,66,40,168),(81,0,0,0),(0,3,0,0),(2,3,0,0),(2,3,143,0),(241,3,143,0),(241,75,143,0),(241,75,246,0),(241,233,246,0),(241,233,246,95),(204,233,246,95),(204,233,246,50),(204,233,20,50),(204,91,20,50),(204,21,20,50),(204,21,113,50),(204,21,113,69),(7,21,113,69),(7,21,113,135),(7,21,113,208),(0,123,0,0),(110,123,0,0),(0,0,0,127),(0,0,0,242),(138,0,0,242),(138,0,107,242),(138,0,107,108),(138,154,107,108),(205,0,0,0),(144,0,0,0),(34,0,0,0),(34,0,143,0),(34,0,191,0),(34,0,191,72),(34,0,191,85),(34,0,191,126),(34,12,191,126),(102,12,191,126),(102,82,191,126),(102,82,191,134),(40,82,191,134),(40,104,191,134),(40,104,191,149),(40,18,191,149),(162,18,191,149),(162,159,191,149),(162,130,191,149),(162,135,191,149),(162,135,25,149),(162,135,25,251),(162,135,173,251),(162,135,100,251),(162,135,100,150),(162,135,182,150),(225,135,182,150),(152,135,182,150),(152,135,182,203),(152,213,182,203),(0,0,0,245),(0,0,0,22),(0,141,0,22),(0,245,0,22),(166,245,0,22),(116,245,0,22),(158,245,0,22),(158,2,0,22),(158,2,59,22),(0,0,2,0),(0,0,71,0),(0,136,71,0),(0,136,200,0),(99,136,200,0),(99,136,197,0),(99,136,98,0),(99,136,145,0),(0,151,0,0),(133,151,0,0),(133,151,0,167),(241,151,0,167),(195,151,0,167),(195,151,0,7),(195,104,0,7),(195,104,193,7),(195,154,193,7),(195,240,193,7),(195,107,193,7),(125,107,193,7),(47,107,193,7),(6,107,193,7),(6,107,30,7),(6,36,30,7),(23,36,30,7),(23,36,30,242),(0,0,0,69),(0,130,0,69),(0,174,0,69),(0,174,0,72),(47,174,0,72),(47,72,0,72),(108,72,0,72),(0,0,200,0),(22,0,200,0),(22,0,200,253),(22,0,181,253),(22,0,181,67),(22,139,181,67),(3,139,181,67),(3,139,181,16),(3,139,49,16),(207,139,49,16),(207,155,49,16),(63,155,49,16),(63,88,49,16),(63,88,10,16),(63,88,10,147),(63,88,181,147),(63,191,181,147),(144,191,181,147),(144,65,181,147),(173,65,181,147),(173,65,11,147),(173,65,205,147),(173,65,205,122),(0,72,0,0),(45,72,0,0),(45,72,0,191),(45,181,0,191),(45,60,0,191),(45,46,0,191),(45,107,0,191),(45,107,84,191),(45,107,173,191),(232,107,173,191),(232,107,173,20),(187,107,173,20),(187,107,24,20),(187,107,103,20),(187,107,55,20),(187,107,238,20),(187,107,238,71),(187,107,238,239),(250,107,238,239),(250,195,238,239),(89,195,238,239),(89,195,144,239),(89,195,144,175),(138,195,144,175),(138,195,66,175),(247,195,66,175),(247,195,66,84),(247,195,66,160),(247,195,66,87),(247,109,66,87),(0,0,140,0),(208,0,140,0),(208,0,140,200),(208,0,217,200),(208,170,217,200),(208,170,217,72),(0,0,0,171),(126,0,0,171),(207,0,0,171),(45,0,0,171),(45,0,0,174),(45,0,0,237),(45,0,0,200),(0,0,0,142),(0,122,0,142),(214,0,0,0),(214,0,0,45),(214,0,75,45),(214,0,75,186),(214,0,75,84),(15,0,75,84),(15,0,62,84),(132,0,62,84),(46,0,62,84),(19,0,62,84),(19,0,133,84),(138,0,133,84),(138,219,133,84),(50,219,133,84),(12,219,133,84),(12,219,133,93),(12,219,133,154),(12,219,225,154),(0,0,0,226),(0,0,89,226),(0,0,89,35),(36,0,89,35),(36,0,115,35),(36,156,115,35),(32,156,115,35),(32,156,115,77),(32,156,246,77),(32,182,246,77),(32,61,246,77),(32,61,238,77),(0,79,0,0),(0,79,0,98),(0,79,0,248),(0,49,0,0),(189,49,0,0),(189,49,222,0),(189,49,171,0),(189,49,171,119),(189,49,69,119),(189,72,69,119),(226,72,69,119),(248,72,69,119),(248,72,69,235),(248,245,69,235),(41,245,69,235),(41,245,69,16),(41,245,69,70),(192,245,69,70),(192,220,69,70),(192,220,69,46),(192,116,69,46),(131,116,69,46),(131,203,69,46),(27,203,69,46),(27,125,69,46),(27,125,69,222),(231,125,69,222),(143,125,69,222),(143,125,69,144),(143,209,69,144),(229,209,69,144),(229,209,69,193),(229,177,69,193),(229,0,0,0),(224,0,0,0),(183,0,0,0),(183,0,239,0),(0,0,93,0),(186,0,93,0),(186,0,93,64),(247,0,93,64),(247,0,84,64),(247,147,84,64),(0,0,181,0),(0,159,181,0),(139,159,181,0),(139,159,181,240),(53,159,181,240),(162,159,181,240),(162,47,181,240),(162,47,203,240),(162,50,203,240),(162,233,203,240),(162,233,124,240),(241,233,124,240),(0,0,0,170),(0,227,0,170),(0,0,0,227),(95,0,0,227),(95,103,0,227),(95,103,0,84),(95,13,0,84),(181,13,0,84),(51,13,0,84),(0,0,0,239),(11,0,0,239),(0,0,0,64),(73,0,0,64),(73,0,0,157),(73,52,0,157),(73,52,0,53),(73,52,0,64),(73,52,51,64),(73,52,51,101),(73,240,51,101),(0,0,0,200),(0,208,0,200),(0,208,14,200),(0,95,14,200),(0,95,165,200),(0,44,165,200),(0,113,165,200),(0,113,165,32),(0,11,165,32),(0,11,165,32),(0,11,242,32),(110,11,242,32),(0,177,0,0),(0,177,0,32),(130,177,0,32),(130,177,0,41),(120,177,0,41),(0,0,0,95),(147,0,0,0),(222,0,0,0),(0,0,146,0),(0,126,146,0),(0,233,146,0),(0,123,146,0),(191,123,146,0),(191,123,223,0),(191,158,223,0),(191,90,223,0),(191,90,223,100),(191,98,223,100),(191,113,223,100),(191,113,223,122),(191,22,223,122),(191,22,186,122),(191,22,186,46),(10,22,186,46),(10,22,186,181),(10,22,186,35),(10,22,79,35),(10,22,79,195),(80,22,79,195),(80,193,79,195),(80,193,81,195),(243,193,81,195),(243,193,81,164),(243,193,101,164),(46,193,101,164),(46,193,240,164),(46,193,223,164),(75,193,223,164),(22,193,223,164),(94,193,223,164),(84,193,223,164),(84,193,14,164),(84,15,14,164),(84,47,14,164),(84,47,204,164),(84,47,204,196),(84,47,102,196),(201,47,102,196),(201,119,102,196),(201,52,102,196),(201,226,102,196),(201,226,102,106),(201,226,162,106),(201,226,162,98),(201,226,162,220),(201,226,115,220),(201,226,115,10),(201,210,115,10),(201,210,154,10),(201,210,154,250),(146,210,154,250),(209,210,154,250),(209,59,154,250),(209,59,154,214),(209,59,154,76),(234,59,154,76),(234,59,221,76),(234,59,79,76),(0,48,0,0),(0,48,38,0),(0,48,14,0),(0,48,14,104),(0,48,122,104),(0,71,122,104),(0,174,122,104),(0,174,122,210),(0,121,122,210),(54,121,122,210),(54,121,137,210),(54,138,137,210),(54,18,137,210),(54,18,137,12),(54,200,137,12),(54,55,137,12),(190,55,137,12),(190,55,199,12),(190,55,199,115),(190,199,199,115),(190,199,199,10),(197,199,199,10),(197,199,137,10),(197,177,137,10),(197,89,137,10),(197,89,74,10),(139,89,74,10),(147,89,74,10),(147,111,74,10),(147,1,74,10),(251,1,74,10),(251,1,74,240),(48,1,74,240),(48,186,74,240),(119,186,74,240),(52,186,74,240),(52,201,74,240),(52,201,74,48),(32,201,74,48),(32,201,119,48),(32,77,119,48),(32,74,119,48),(32,143,119,48),(201,0,0,0),(201,0,0,237),(201,0,45,237),(201,0,36,237),(201,0,36,40),(201,0,21,40),(201,0,21,227),(201,186,21,227),(201,186,48,227),(201,21,48,227),(0,0,170,0),(0,0,170,4),(0,201,170,4),(0,149,170,4),(105,149,170,4),(0,0,135,0),(0,0,135,155),(0,0,238,155),(0,0,215,155),(0,216,215,155),(0,216,208,155),(0,216,208,113),(222,216,208,113),(222,216,208,109),(0,0,14,0),(0,0,14,75),(0,0,138,75),(144,0,138,75),(144,156,138,75),(78,156,138,75),(78,156,138,100),(0,0,64,0),(112,0,64,0),(112,0,64,91),(112,82,64,91),(0,0,0,14),(0,43,0,14),(0,43,117,14),(0,232,117,14),(0,232,155,14),(0,232,155,47),(0,0,0,73),(0,0,0,243),(0,102,0,243),(212,102,0,243),(239,102,0,243),(239,102,254,243),(0,0,19,0),(0,189,19,0),(0,189,19,102),(0,189,19,133),(0,135,19,133),(0,135,190,133),(0,135,67,133),(0,146,67,133),(0,146,67,233),(0,146,67,54),(0,146,67,118),(0,146,218,118),(0,146,218,95),(30,146,218,95),(111,146,218,95),(111,146,203,95),(0,30,0,0),(0,239,0,0),(0,0,0,69),(0,0,196,0),(0,8,196,0),(0,8,135,0),(0,8,1,0),(0,8,1,48),(0,213,1,48),(0,147,1,48),(0,147,1,71),(0,147,255,71),(0,147,24,71),(0,147,24,145),(0,147,63,145),(0,0,58,0),(98,0,58,0),(98,0,235,0),(98,0,149,0),(98,48,149,0),(98,48,230,0),(0,0,0,2),(0,45,0,2),(0,239,0,2),(159,239,0,2),(34,239,0,2),(194,239,0,2),(238,239,0,2),(238,239,111,2),(238,239,111,190),(238,239,111,196),(238,239,72,196),(132,239,72,196),(132,0,72,196),(43,0,72,196),(43,0,137,196),(119,0,137,196),(119,0,137,199),(232,0,137,199),(232,0,197,199),(253,0,197,199),(189,0,197,199),(189,0,197,114),(189,0,197,4),(189,0,197,237),(189,218,197,237),(189,218,172,237),(189,228,172,237),(6,228,172,237),(6,228,172,144),(6,60,172,144),(59,60,172,144),(59,60,172,18),(48,60,172,18),(0,140,0,0),(0,140,0,181),(0,140,0,252),(0,11,0,252),(146,11,0,252),(146,11,0,228),(146,11,0,26),(146,11,0,13),(146,12,0,13),(146,12,30,13),(146,135,30,13),(146,135,169,13),(146,135,166,13),(146,249,166,13),(188,249,166,13),(75,249,166,13),(75,249,166,108),(32,249,166,108),(32,249,153,108),(32,249,168,108),(249,249,168,108),(249,173,168,108),(12,173,168,108),(12,93,168,108),(12,93,168,188),(12,93,111,188),(12,93,189,188),(12,199,189,188),(12,199,195,188),(12,199,238,188),(12,199,238,246),(12,199,238,141),(12,165,238,141),(12,6,238,141),(12,6,238,3),(12,6,125,3),(12,6,118,3),(12,6,118,69),(12,219,118,69),(12,219,36,69),(12,219,43,69),(12,219,43,5),(225,219,43,5),(225,219,54,5),(201,219,54,5),(51,219,54,5),(51,219,54,36),(217,219,54,36),(231,219,54,36),(0,0,0,159),(0,0,226,159),(0,0,0,159),(0,0,217,159),(0,170,217,159),(0,170,217,6),(0,170,217,30),(0,170,141,30),(0,170,141,235),(0,170,104,235),(0,209,104,235),(41,0,0,0),(41,0,0,113),(121,0,0,113),(121,0,0,247),(58,0,0,247),(58,87,0,247),(58,87,0,149),(58,10,0,149),(143,10,0,149),(143,51,0,149),(143,51,44,149),(84,51,44,149),(84,150,44,149),(84,150,44,238),(84,254,44,238),(84,227,44,238),(0,0,0,126),(0,196,0,126),(0,196,0,159),(0,196,32,159),(204,196,32,159),(33,196,32,159),(151,196,32,159),(151,16,32,159),(151,16,32,171),(151,94,32,171),(243,94,32,171),(243,94,32,37),(0,0,125,0),(0,0,0,146),(125,0,0,146),(125,0,167,146),(143,0,167,146),(143,23,167,146),(63,23,167,146),(63,23,167,39),(63,23,85,39),(54,0,0,0),(54,6,0,0),(54,6,28,0),(135,6,28,0),(135,6,64,0),(135,6,64,183),(0,160,0,0),(0,160,191,0),(0,122,191,0),(0,122,134,0),(0,122,197,0),(0,122,197,206),(157,122,197,206),(157,122,40,206),(157,221,40,206),(157,221,40,242),(157,221,58,242),(217,221,58,242),(0,0,0,9),(0,0,235,9),(0,0,7,9),(0,0,7,254),(104,0,7,254),(219,0,7,254),(219,0,7,237),(219,0,165,237),(219,0,226,237),(219,0,138,237),(219,0,138,237),(198,0,0,0),(100,0,0,0),(100,0,0,159),(100,0,0,185),(15,0,0,185),(15,173,0,185),(112,173,0,185),(1,0,0,0),(1,102,0,0),(1,210,0,0),(0,0,3,0),(0,160,3,0),(54,160,3,0),(54,160,3,12),(54,160,31,12),(0,0,0,2),(0,0,0,66),(0,140,0,66),(119,140,0,66),(0,0,245,0),(0,8,245,0),(9,8,245,0),(9,8,245,254),(9,8,95,254),(9,8,95,245),(3,8,95,245),(3,8,95,239),(3,108,95,239),(3,108,95,194),(81,108,95,194),(81,108,95,163),(81,189,95,163),(81,189,95,188),(18,189,95,188),(18,13,95,188),(18,13,95,120),(27,13,95,120),(27,13,95,212),(70,13,95,212),(12,13,95,212),(32,13,95,212),(0,0,226,0),(4,0,226,0),(4,190,226,0),(0,16,0,0),(0,84,0,0),(51,84,0,0),(51,26,0,0),(190,26,0,0),(190,26,0,175),(0,13,0,0),(0,13,214,0),(0,200,214,0),(0,200,191,0),(0,169,191,0),(0,179,191,0),(107,179,191,0),(28,179,191,0),(0,0,154,0),(50,0,154,0),(50,0,154,92),(50,0,154,48),(198,0,154,48),(198,0,199,48),(198,0,13,48),(198,0,13,115),(198,126,13,115),(198,84,13,115),(198,55,13,115),(198,55,13,105),(198,55,175,105),(198,55,73,105),(185,55,73,105),(185,36,73,105),(204,36,73,105),(117,36,73,105),(117,70,73,105),(117,83,73,105),(117,83,255,105),(117,83,255,202),(117,129,255,202),(197,129,255,202),(197,129,255,57),(197,129,255,161),(197,49,255,161),(197,49,13,161),(0,74,0,0),(0,74,0,17),(0,74,59,17),(0,74,59,36),(0,74,59,205),(0,74,59,159),(0,74,211,159),(0,167,211,159),(0,167,211,189),(0,167,181,189),(0,167,181,220),(117,167,181,220),(144,167,181,220),(144,163,181,220),(144,163,181,10),(217,163,181,10),(0,0,181,0),(0,0,25,0),(227,0,25,0),(56,0,25,0),(234,0,25,0),(234,0,25,22),(234,0,25,194),(234,208,25,194),(234,208,25,32),(234,131,25,32),(234,131,201,32),(234,131,191,32),(194,131,191,32),(194,131,191,124),(194,131,114,124),(194,131,114,14),(194,131,225,14),(194,131,225,101),(194,131,121,101),(194,131,121,196),(91,131,121,196),(180,131,121,196),(180,131,121,243),(180,131,121,128),(0,0,229,0),(0,0,33,0),(0,0,10,0),(0,0,10,49),(0,0,10,95),(0,0,10,21),(99,0,10,21),(170,0,10,21),(170,64,10,21),(170,64,10,143),(170,64,64,143),(170,64,64,42),(170,64,64,52),(170,64,64,10),(137,64,64,10),(210,64,64,10),(210,64,64,127),(210,102,64,127),(210,193,64,127),(210,188,64,127),(210,188,223,127),(64,188,223,127),(64,188,246,127),(64,188,246,25),(206,188,246,25),(75,188,246,25),(75,180,246,25),(75,107,246,25),(75,27,246,25),(0,0,0,143),(0,0,44,0),(0,0,250,0),(199,0,250,0),(199,0,250,138),(199,0,250,243),(199,0,228,243),(199,0,228,205),(199,0,228,173),(0,0,249,0),(0,0,55,0),(0,0,78,0),(156,0,78,0),(156,0,78,224),(156,0,78,76),(0,0,0,128),(0,0,208,128),(0,0,246,128),(0,162,246,128),(0,164,246,128),(0,164,246,113),(0,164,246,231),(0,164,157,231),(0,0,0,181),(0,99,0,181),(0,12,0,181),(93,12,0,181),(163,12,0,181),(163,12,95,181),(163,46,95,181),(61,0,0,0),(61,145,0,0),(225,145,0,0),(225,247,0,0),(225,245,0,0),(225,245,0,98),(225,245,149,98),(225,245,252,98),(225,245,26,98),(0,0,0,152),(0,0,0,69),(0,228,0,69),(0,164,0,69),(198,164,0,69),(198,164,0,58),(198,232,0,58),(198,101,0,58),(198,101,160,58),(198,218,160,58),(147,218,160,58),(53,218,160,58),(53,218,160,37),(53,104,160,37),(53,236,160,37),(0,0,89,0),(235,0,0,0),(0,0,0,74),(0,0,0,122),(0,0,0,93),(234,0,0,93),(234,0,0,120),(234,251,0,120),(234,251,169,120),(234,230,169,120),(234,198,169,120),(234,198,169,8),(234,129,169,8),(234,129,169,240),(234,129,169,216),(86,129,169,216),(86,54,169,216),(0,0,0,157),(128,0,0,157),(128,0,229,157),(200,0,229,157),(200,0,229,31),(36,0,0,0),(48,0,0,0),(243,0,0,0),(243,41,0,0),(0,154,0,0),(0,103,0,0),(0,103,0,37),(0,131,0,37),(0,224,0,37),(0,0,190,0),(0,0,190,120),(0,210,190,120),(0,210,221,120),(66,210,221,120),(66,45,221,120),(66,253,221,120),(174,253,221,120),(174,200,221,120),(246,200,221,120),(246,2,221,120),(246,2,221,247),(246,2,118,247),(246,2,146,247),(237,2,146,247),(55,2,146,247),(55,2,243,247),(55,2,243,40),(55,2,202,40),(55,2,88,40),(55,2,88,123),(252,2,88,123),(205,2,88,123),(205,117,88,123),(139,117,88,123),(139,0,88,123),(28,0,88,123),(138,0,88,123),(151,0,88,123),(0,0,0,135),(0,0,75,135),(0,151,75,135),(0,40,75,135),(0,40,216,135),(0,40,216,193),(0,40,216,82),(0,40,216,55),(0,86,216,55),(0,66,216,55),(0,66,109,55),(0,66,58,55),(0,66,58,218),(0,60,58,218),(0,79,58,218),(0,35,58,218),(228,35,58,218),(243,35,58,218),(243,35,16,218),(243,35,16,215),(243,35,250,215),(243,193,250,215),(243,193,213,215),(243,140,213,215),(243,140,207,215),(19,140,207,215),(19,140,47,215),(19,140,47,19),(19,140,47,233),(0,143,0,0),(25,143,0,0),(25,143,0,3),(0,132,0,0),(248,132,0,0),(248,132,0,188),(152,132,0,188),(252,132,0,188),(252,178,0,188),(69,178,0,188),(69,45,0,188),(69,45,103,188),(69,45,228,188),(69,45,64,188),(167,45,64,188),(200,45,64,188),(200,252,64,188),(205,0,0,0),(205,88,0,0),(205,88,0,31),(55,88,0,31),(229,88,0,31),(249,88,0,31),(0,88,0,31),(0,88,152,31),(87,88,152,31),(87,5,152,31),(0,0,0,251),(0,0,182,251),(67,0,182,251),(67,0,182,169),(67,229,182,169),(67,229,182,195),(242,229,182,195),(242,250,182,195),(242,225,182,195),(5,225,182,195),(245,0,0,0),(245,220,0,0),(245,220,0,209),(211,220,0,209),(211,220,237,209),(211,220,62,209),(10,220,62,209),(64,220,62,209),(64,220,62,70),(64,220,62,228),(64,220,62,152),(206,220,62,152),(206,220,139,152),(75,220,139,152),(0,0,0,87),(0,31,0,87),(0,180,0,87),(0,180,0,186),(73,180,0,186),(73,180,0,121),(170,180,0,121),(170,180,143,121),(170,247,143,121),(170,247,143,226),(170,250,143,226),(170,41,143,226),(170,41,143,168),(170,177,143,168),(170,177,133,168),(170,87,133,168),(170,87,133,249),(170,87,39,249),(170,87,2,249),(170,87,127,249),(170,97,127,249),(165,97,127,249),(165,97,103,249),(168,97,103,249),(168,136,103,249),(168,136,103,144),(124,136,103,144),(124,144,103,144),(124,119,103,144),(124,34,103,144),(124,126,103,144),(124,126,252,144),(124,58,252,144),(124,58,204,144),(31,58,204,144),(31,181,204,144),(31,181,15,144),(228,181,15,144),(228,181,195,144),(10,181,195,144),(10,181,195,46),(10,181,195,46),(10,73,195,46),(10,73,254,46),(10,73,130,46),(10,73,130,87),(10,73,34,87),(10,73,108,87),(10,73,43,87),(42,73,43,87),(42,211,43,87),(231,211,43,87),(231,211,120,87),(0,117,0,0),(0,117,34,0),(0,117,47,0),(0,117,47,19),(0,230,0,0),(0,230,51,0),(0,230,51,248),(0,230,3,248),(0,230,3,13),(0,230,3,116),(0,230,240,116),(0,230,240,2),(0,230,197,2),(83,230,197,2),(123,230,197,2),(123,20,197,2),(123,20,233,2),(244,20,233,2),(244,20,162,2),(69,20,162,2),(69,20,210,2),(69,20,210,117),(207,20,210,117),(237,20,210,117),(125,20,210,117),(125,239,210,117),(125,117,210,117),(36,0,0,0),(36,0,229,0),(36,0,5,0),(36,0,75,0),(36,0,153,0),(36,170,153,0),(0,0,40,0),(0,0,92,0),(0,0,92,255),(0,130,92,255),(0,130,29,255),(135,130,29,255),(135,130,210,255),(135,130,210,93),(135,125,210,93),(39,125,210,93),(82,125,210,93),(82,125,210,241),(82,125,79,241),(82,213,79,241),(60,213,79,241),(60,213,8,241),(60,242,8,241),(60,242,206,241),(60,242,122,241),(60,242,122,116),(0,0,87,0),(0,0,87,145),(0,183,87,145),(0,183,14,145),(37,183,14,145),(223,183,14,145),(245,183,14,145),(245,183,197,145),(5,183,197,145),(150,183,197,145),(150,105,197,145),(239,105,197,145),(239,27,197,145),(239,145,197,145),(239,145,70,145),(239,177,70,145),(239,177,161,145),(239,177,188,145),(88,177,188,145),(88,177,188,199),(88,177,188,5),(88,177,185,5),(88,81,185,5),(88,81,248,5),(122,81,248,5),(122,81,204,5),(0,0,0,249),(145,0,0,249),(246,0,0,249),(246,218,0,249),(134,218,0,249),(70,0,0,0),(178,0,0,0),(178,254,0,0),(164,254,0,0),(164,254,0,198),(164,254,0,7),(172,254,0,7),(172,254,130,7),(172,57,130,7),(172,67,130,7),(5,67,130,7),(5,67,130,157),(5,67,34,157),(26,67,34,157),(26,67,36,157),(26,67,59,157),(131,67,59,157),(131,163,59,157),(131,163,59,158),(100,163,59,158),(100,218,59,158),(220,218,59,158),(244,218,59,158),(244,218,59,39),(244,32,59,39),(102,32,59,39),(102,32,231,39),(102,32,231,192),(230,32,231,192),(210,32,231,192),(9,32,231,192),(18,32,231,192),(18,32,231,80),(18,32,145,80),(18,32,161,80),(18,32,54,80),(18,32,155,80),(18,32,107,80),(18,32,34,80),(18,32,45,80),(18,240,45,80),(18,240,207,80),(18,240,242,80),(18,240,241,80),(18,240,241,46),(49,240,241,46),(49,240,241,45),(152,240,241,45),(152,240,241,92),(152,249,241,92),(198,249,241,92),(198,249,241,241),(198,68,241,241),(244,0,0,0),(28,0,0,0),(28,0,174,0),(28,0,174,120),(39,0,174,120),(39,0,174,121),(181,0,174,121),(218,0,174,121),(218,127,174,121),(66,127,174,121),(66,127,20,121),(66,127,232,121),(0,0,0,245),(0,0,208,245),(0,122,208,245),(143,122,208,245),(143,122,224,245),(143,10,224,245),(143,149,224,245),(143,149,101,245),(143,149,101,54),(26,149,101,54),(123,149,101,54),(123,149,101,95),(28,149,101,95),(195,149,101,95),(195,149,101,126),(119,149,101,126),(119,149,101,221),(119,149,101,84),(0,0,253,0),(0,0,253,170),(0,0,125,170),(0,0,230,170),(0,0,0,186),(0,231,0,186),(170,231,0,186),(170,107,0,186),(170,107,190,186),(170,108,190,186),(170,108,224,186),(170,188,224,186),(108,188,224,186),(108,232,224,186),(108,212,224,186),(240,212,224,186),(240,212,224,202),(252,212,224,202),(252,212,163,202),(252,212,163,94),(252,212,163,5),(65,212,163,5),(50,212,163,5),(50,126,163,5),(0,131,0,0),(0,176,0,0),(0,176,153,0),(0,176,153,78),(0,173,153,78),(0,0,78,0),(0,0,17,0),(0,0,224,0),(218,0,224,0),(218,16,224,0),(94,16,224,0),(94,236,224,0),(152,236,224,0),(152,232,224,0),(152,7,224,0),(152,123,224,0),(86,123,224,0),(86,123,224,109),(176,123,224,109),(176,123,224,90),(34,123,224,90),(34,123,152,90),(23,123,152,90),(77,123,152,90),(77,123,21,90),(77,114,21,90),(77,20,21,90),(77,20,21,214),(77,20,21,34),(77,190,21,34),(77,190,116,34),(243,190,116,34),(243,190,116,197),(0,83,0,0),(0,83,0,138),(0,146,0,0),(0,146,8,0),(0,146,8,152),(172,146,8,152),(208,146,8,152),(5,146,8,152),(5,194,8,152),(5,194,211,152),(5,231,211,152),(159,231,211,152),(159,231,211,196),(249,231,211,196),(0,0,194,0),(0,59,194,0),(0,137,194,0),(0,137,226,0),(0,137,226,61),(0,137,226,48),(0,15,226,48),(0,15,237,48),(39,0,0,0),(39,0,228,0),(39,0,190,0),(0,0,0,178),(0,216,0,178),(0,216,28,178),(0,216,199,178),(169,216,199,178),(236,216,199,178),(236,78,199,178),(236,77,199,178),(236,77,199,49),(190,77,199,49),(58,77,199,49),(58,77,199,200),(58,225,199,200),(7,225,199,200),(7,225,213,200),(22,225,213,200),(234,225,213,200),(234,225,1,200),(0,111,0,0),(0,111,0,9),(0,116,0,9),(0,116,185,9),(0,116,195,9),(0,116,195,203),(0,116,195,117),(0,116,53,117),(0,116,53,26),(0,116,221,26),(0,204,221,26),(0,40,221,26),(0,40,227,26),(39,40,227,26),(39,194,227,26),(0,126,0,0),(0,181,0,0),(0,181,210,0),(0,181,150,0),(137,181,150,0),(137,181,192,0),(137,181,192,189),(159,181,192,189),(159,181,192,159),(159,181,192,3),(14,181,192,3),(14,247,192,3),(42,247,192,3),(0,0,105,0),(221,0,105,0),(221,0,31,0),(221,0,102,0),(221,0,167,0),(221,107,167,0),(221,107,167,93),(221,107,167,135),(180,107,167,135),(180,107,167,139),(180,107,131,139),(178,107,131,139),(178,107,93,139),(162,107,93,139),(94,107,93,139),(94,107,93,60),(209,107,93,60),(209,107,189,60),(209,107,189,93),(209,107,7,93),(209,76,7,93),(121,76,7,93),(121,76,227,93),(121,76,227,76),(121,76,227,68),(121,76,227,63),(163,76,227,63),(163,76,16,63),(221,76,16,63),(221,76,159,63),(221,72,159,63),(54,0,0,0),(54,0,106,0),(54,0,110,0),(0,0,5,0),(0,97,5,0),(0,97,227,0),(0,97,227,206),(164,97,227,206),(164,97,227,114),(164,97,227,94),(164,97,208,94),(164,97,251,94),(164,97,192,94),(164,97,192,5),(146,97,192,5),(146,200,192,5),(146,200,128,5),(146,200,128,220),(146,200,102,220),(149,200,102,220),(149,200,28,220),(149,200,156,220),(149,200,22,220),(149,200,44,220),(127,200,44,220),(127,200,44,99),(88,0,0,0),(128,0,0,0),(128,0,0,122),(128,50,0,122),(128,50,91,122),(128,50,224,122),(128,50,253,122),(0,232,0,0),(0,186,0,0),(0,227,0,0),(0,227,0,169),(0,214,0,169),(79,214,0,169),(79,190,0,169),(79,190,0,137),(79,190,206,137),(54,190,206,137),(114,190,206,137),(114,190,123,137),(114,247,123,137),(114,247,151,137),(0,157,0,0),(0,157,0,95),(0,157,123,95),(0,216,123,95),(0,216,123,30),(185,216,123,30),(172,216,123,30),(172,63,123,30),(172,63,123,78),(125,63,123,78),(125,63,169,78),(242,63,169,78),(242,63,169,135),(242,115,169,135),(242,115,45,135),(242,115,45,221),(242,238,45,221),(242,238,62,221),(242,238,34,221),(242,150,34,221),(242,57,34,221),(16,57,34,221),(16,18,34,221),(16,18,34,23),(16,18,132,23),(16,83,132,23),(122,83,132,23),(122,52,132,23),(30,52,132,23),(62,52,132,23),(62,52,132,201),(62,52,132,201),(62,103,132,201),(110,103,132,201),(110,103,112,201),(110,103,203,201),(110,103,238,201),(110,120,238,201),(110,120,238,186),(110,120,210,186),(110,120,30,186),(0,171,0,0),(0,171,0,166),(0,221,0,166),(0,221,0,237),(0,202,0,237),(166,202,0,237),(166,120,0,237),(166,120,0,179),(156,120,0,179),(156,120,0,105),(156,120,0,124),(156,120,0,124),(156,120,0,65),(17,120,0,65),(17,143,0,65),(17,143,30,65),(17,143,45,65),(17,243,45,65),(17,243,45,209),(17,172,45,209),(0,0,0,125),(0,0,0,240),(0,80,0,0),(205,80,0,0),(205,80,0,11),(205,232,0,11),(10,232,0,11),(0,0,0,4),(0,0,55,4),(0,0,55,117),(0,0,30,117),(178,0,30,117),(178,0,73,117),(178,47,73,117),(178,47,90,117),(178,70,90,117),(178,70,133,117),(178,202,133,117),(178,202,129,117),(178,202,129,156),(253,202,129,156),(253,202,129,237),(253,202,83,237),(253,179,83,237),(93,179,83,237),(93,15,83,237),(11,0,0,0),(0,0,106,0),(0,0,182,0),(83,0,182,0),(83,64,182,0),(83,64,182,87),(83,64,182,60),(83,64,144,60),(83,64,54,60),(83,64,54,225),(125,64,54,225),(125,213,54,225),(125,180,54,225),(125,180,5,225),(125,180,163,225),(125,180,245,225),(136,180,245,225),(136,180,89,225),(212,180,89,225),(212,180,178,225),(212,180,18,225),(212,180,148,225),(212,2,148,225),(217,2,148,225),(217,2,148,250),(217,204,148,250),(217,204,77,250),(143,204,77,250),(160,204,77,250),(160,204,77,53),(0,0,0,75),(0,0,0,133),(0,0,0,151),(0,0,182,151),(255,0,0,0),(255,0,0,139),(255,0,0,206),(50,0,0,206),(50,0,230,206),(50,223,230,206),(50,23,230,206),(50,221,230,206),(48,221,230,206),(48,221,230,92),(48,71,230,92),(0,82,0,0),(0,0,34,0),(0,0,34,31),(0,0,27,31),(0,0,27,127),(0,0,27,208),(50,0,27,208),(50,47,27,208),(209,47,27,208),(209,47,27,11),(209,47,27,162),(39,47,27,162),(39,47,27,62),(39,47,27,29),(39,207,27,29),(39,207,14,29),(39,207,92,29),(39,207,92,18),(39,207,92,192),(39,207,107,192),(39,207,157,192),(75,207,157,192),(75,207,157,167),(75,207,180,167),(148,207,180,167),(148,79,180,167),(148,79,180,89),(148,79,180,140),(148,79,180,5),(148,79,180,239),(148,138,180,239),(148,138,196,239),(0,104,0,0),(172,104,0,0),(172,104,0,89),(172,104,0,207),(172,104,0,77),(172,7,0,77),(172,7,130,77),(0,0,106,0),(0,151,106,0),(168,151,106,0),(233,151,106,0),(76,151,106,0),(76,151,65,0),(213,151,65,0),(213,151,65,139),(213,151,147,139),(162,151,147,139),(44,151,147,139),(202,151,147,139),(202,112,147,139),(202,112,147,216),(83,112,147,216),(47,112,147,216),(43,112,147,216),(43,3,147,216),(43,3,147,161),(43,3,114,161),(43,3,76,161),(43,3,76,41),(43,3,76,85),(43,58,76,85),(0,0,0,51),(0,0,0,63),(0,0,93,63),(65,0,93,63),(65,250,93,63),(103,250,93,63),(48,250,93,63),(48,250,10,63),(175,250,10,63),(175,250,10,246),(137,250,10,246),(137,250,10,223),(137,250,64,223),(0,0,199,0),(0,196,199,0),(201,196,199,0),(201,196,88,0),(201,196,88,236),(201,196,210,236),(0,0,0,54),(0,0,0,77),(0,0,196,0),(0,181,196,0),(0,78,0,0),(0,78,22,0),(0,78,41,0),(175,78,41,0),(175,78,41,221),(175,105,41,221),(175,105,85,221),(175,196,85,221),(175,196,181,221),(56,196,181,221),(224,196,181,221),(224,196,40,221),(224,196,40,4),(207,0,0,0),(207,25,0,0),(207,25,173,0),(207,25,173,163),(207,25,34,163),(207,250,34,163),(0,47,0,0),(0,218,0,0),(92,218,0,0),(92,218,0,80),(92,218,0,158),(92,218,0,223),(92,218,16,223),(0,0,0,80),(0,0,0,126),(135,0,0,126),(135,0,176,126),(135,0,176,185),(0,96,0,0),(0,96,48,0),(0,251,0,0),(0,131,0,0),(0,131,88,0),(0,131,88,8),(50,131,88,8),(27,131,88,8),(27,131,100,8),(27,131,13,8),(27,131,101,8),(27,166,101,8),(46,166,101,8),(188,166,101,8),(188,166,101,75),(188,63,101,75),(188,63,101,195),(91,63,101,195),(91,63,137,195),(91,63,57,195),(91,199,57,195),(155,199,57,195),(155,218,57,195),(221,218,57,195),(221,218,57,69),(221,26,57,69),(221,103,57,69),(221,103,57,112),(238,103,57,112),(238,103,123,112),(238,103,123,188),(238,103,223,188),(238,47,223,188),(238,139,223,188),(149,139,223,188),(149,139,223,234),(240,139,223,234),(240,139,206,234),(240,139,206,235),(240,139,147,235),(240,139,219,235),(240,142,219,235),(240,142,74,235),(240,142,74,33),(187,142,74,33),(211,142,74,33),(211,142,74,232),(0,198,0,0),(181,198,0,0),(181,159,0,0),(154,159,0,0),(154,159,183,0),(154,159,197,0),(154,118,197,0),(0,0,60,0),(0,0,60,68),(0,0,251,68),(162,0,251,68),(162,0,251,157),(20,0,251,157),(20,225,251,157),(20,225,64,157),(20,225,64,238),(173,225,64,238),(173,225,18,238),(111,225,18,238),(111,225,18,90),(111,187,18,90),(111,32,18,90),(111,32,90,90),(148,32,90,90),(73,32,90,90),(0,0,0,230),(0,0,91,230),(0,0,175,230),(150,0,175,230),(150,0,175,127),(30,0,175,127),(194,0,175,127),(218,0,175,127),(142,0,175,127),(142,0,175,18),(142,0,175,11),(142,0,241,11),(142,97,241,11),(142,181,241,11),(142,181,235,11),(142,88,235,11),(8,88,235,11),(169,88,235,11),(169,123,235,11),(169,155,235,11),(169,155,198,11),(169,155,187,11),(169,155,116,11),(169,155,116,31),(169,155,116,31),(169,155,136,31),(169,155,136,114),(169,155,75,114),(169,155,98,114),(169,47,98,114),(0,194,0,0),(0,46,0,0),(46,46,0,0),(46,46,136,0),(194,46,136,0),(194,46,26,0),(82,0,0,0),(158,0,0,0),(158,0,207,0),(203,0,207,0),(203,249,207,0),(153,249,207,0),(153,223,207,0),(153,160,207,0),(153,16,207,0),(0,0,182,0),(0,0,182,237),(0,0,1,237),(57,0,1,237),(57,0,198,237),(0,0,155,0),(0,0,155,185),(224,0,155,185),(224,0,155,87),(53,0,155,87),(53,0,209,87),(53,0,209,181),(53,0,209,38),(53,0,195,38),(53,23,195,38),(53,221,195,38),(0,0,9,0),(0,0,22,0),(0,0,185,0),(0,202,185,0),(0,202,113,0),(0,202,113,11),(71,0,0,0),(71,160,0,0),(71,160,0,133),(71,160,102,133),(71,160,133,133),(71,160,133,255),(71,188,133,255),(226,188,133,255),(226,188,105,255),(226,188,105,173),(226,188,105,171),(160,188,105,171),(160,188,105,202),(160,241,105,202),(160,70,105,202),(160,70,135,202),(160,246,135,202),(37,246,135,202),(5,246,135,202),(5,246,116,202),(5,246,116,160),(5,246,194,160),(5,205,194,160),(5,107,194,160),(139,107,194,160),(139,34,194,160),(139,141,194,160),(139,112,194,160),(139,112,186,160),(139,236,186,160),(139,18,186,160),(139,18,44,160),(95,18,44,160),(95,225,44,160),(95,225,245,160),(28,225,245,160),(61,225,245,160),(61,225,25,160),(191,225,25,160),(165,225,25,160),(165,214,25,160),(0,0,0,106),(111,0,0,106),(111,0,0,12),(111,93,0,12),(86,93,0,12),(86,93,32,12),(147,93,32,12),(147,93,239,12),(147,93,239,6),(147,93,199,6),(147,93,0,6),(0,218,0,0),(0,218,196,0),(0,0,25,0),(0,226,25,0),(0,226,236,0),(106,226,236,0),(62,226,236,0),(0,0,0,146),(0,0,146,146),(64,0,146,146),(64,0,100,146),(64,0,100,77),(172,0,100,77),(233,0,100,77),(233,0,205,77),(140,0,205,77),(140,0,104,77),(193,0,104,77),(193,255,104,77),(193,255,227,77),(193,255,227,232),(193,174,227,232),(193,45,227,232),(193,104,227,232),(193,104,241,232),(193,104,241,89),(12,104,241,89),(12,235,241,89),(7,235,241,89),(7,235,214,89),(0,0,0,73),(0,0,164,73),(9,0,164,73),(9,218,164,73),(9,57,164,73),(81,57,164,73),(81,57,234,73),(208,57,234,73),(208,57,106,73),(208,57,134,73),(167,57,134,73),(167,57,45,73),(167,118,45,73),(236,118,45,73),(236,243,45,73),(174,243,45,73),(174,234,45,73),(174,234,214,73),(174,234,210,73),(56,234,210,73),(56,234,210,127),(56,234,210,210),(206,234,210,210),(206,234,93,210),(159,234,93,210),(159,234,93,116),(159,234,221,116),(252,234,221,116),(127,0,0,0),(127,0,144,0),(127,0,144,81),(127,3,144,81),(28,3,144,81),(103,3,144,81),(103,42,144,81),(103,42,144,235),(103,42,97,235),(173,42,97,235),(36,42,97,235),(201,42,97,235),(201,42,97,253),(201,42,18,253),(201,125,18,253),(201,234,18,253),(201,234,22,253),(201,1,22,253),(0,163,0,0),(0,24,0,0),(66,24,0,0),(66,24,0,230),(152,24,0,230),(152,24,0,246),(152,24,0,197),(152,24,33,197),(152,24,178,197),(152,24,178,30),(152,24,29,30),(152,24,29,205),(207,0,0,0),(207,206,0,0),(207,85,0,0),(207,85,0,184),(207,142,0,184),(207,210,0,184),(207,59,0,184),(129,0,0,0),(129,222,0,0),(129,222,0,0),(129,222,215,0),(4,222,215,0),(126,222,215,0),(126,222,255,0),(126,222,254,0),(143,222,254,0),(143,24,254,0),(143,236,254,0),(143,236,252,0),(143,236,26,0),(143,236,221,0),(143,236,221,41),(136,236,221,41),(136,236,176,41),(136,236,176,212),(136,236,123,212),(136,135,123,212),(136,84,123,212),(136,84,123,92),(136,84,100,92),(136,247,100,92),(136,247,100,13),(136,15,100,13),(136,147,100,13),(136,147,231,13),(136,38,231,13),(203,38,231,13),(203,164,231,13),(233,164,231,13),(163,164,231,13),(163,164,91,13),(163,149,91,13),(163,149,91,91),(163,149,179,91),(26,149,179,91),(26,149,179,187),(26,75,179,187),(0,46,0,0),(0,46,82,0),(0,114,82,0),(0,114,82,82),(0,114,82,200),(0,114,54,200),(0,114,54,142),(184,114,54,142),(249,114,54,142),(249,246,54,142),(168,246,54,142),(168,246,54,34),(168,246,16,34),(168,244,16,34),(168,244,238,34),(48,244,238,34),(183,244,238,34),(232,244,238,34),(251,244,238,34),(251,244,164,34),(197,244,164,34),(197,244,164,102),(197,244,51,102),(16,0,0,0),(16,0,183,0),(16,3,183,0),(0,0,0,0),(0,108,0,0),(0,108,224,0),(0,107,224,0),(0,107,224,243),(0,136,224,243),(115,136,224,243),(115,117,224,243),(115,117,224,242),(115,130,224,242),(70,130,224,242),(70,130,23,242),(70,130,23,19),(11,130,23,19),(94,130,23,19),(215,130,23,19),(215,220,23,19),(163,220,23,19),(163,220,23,74),(163,220,23,69),(163,220,23,180),(127,220,23,180),(127,118,23,180),(127,1,23,180),(127,22,23,180),(127,22,136,180),(208,22,136,180),(208,22,120,180),(242,22,120,180),(102,22,120,180),(118,22,120,180),(118,211,120,180),(118,218,120,180),(209,218,120,180),(209,218,120,230),(26,218,120,230),(142,218,120,230),(142,170,120,230),(252,170,120,230),(200,170,120,230),(167,170,120,230),(160,170,120,230),(227,170,120,230),(227,231,120,230),(0,0,98,0),(0,0,229,0),(162,0,229,0),(162,152,229,0),(162,152,229,101),(162,152,229,135),(0,0,7,0),(0,52,0,0),(0,52,71,0),(0,52,71,84),(247,52,71,84),(247,52,71,213),(247,52,71,157),(195,52,71,157),(95,52,71,157),(95,52,116,157),(95,52,199,157),(95,52,199,76),(95,209,199,76),(102,209,199,76),(0,220,0,0),(0,47,0,0),(0,47,255,0),(0,171,255,0),(0,48,255,0),(0,45,255,0),(0,45,38,0),(0,193,38,0),(134,193,38,0),(134,9,38,0),(134,9,174,0),(209,9,174,0),(209,9,174,175),(31,9,174,175),(31,9,174,29),(102,9,174,29),(0,225,0,0),(0,86,0,0),(0,146,0,0),(0,146,0,81),(0,146,60,81),(0,146,234,81),(0,146,234,181),(152,146,234,181),(0,0,0,96),(0,193,0,96),(0,0,0,158),(23,0,0,158),(23,125,0,158),(23,125,17,158),(0,0,0,33),(0,0,0,35),(0,0,0,9),(0,0,8,9),(3,0,8,9),(3,0,8,135),(3,0,24,135),(0,0,24,135),(10,0,24,135),(10,129,24,135),(10,129,1,135),(10,129,19,135),(50,129,19,135),(50,204,19,135),(50,204,194,135),(50,204,194,161),(50,204,238,161),(31,204,238,161),(31,204,238,52),(221,0,0,0),(221,0,0,242),(213,0,0,242),(72,0,0,242),(72,0,24,242),(72,176,24,242),(162,176,24,242),(122,176,24,242),(122,176,241,242),(122,67,241,242),(122,67,241,86),(122,67,132,86),(122,125,132,86),(122,125,132,184),(122,63,132,184),(122,52,132,184),(122,127,132,184),(110,127,132,184),(92,127,132,184),(92,127,165,184),(92,150,165,184),(92,160,165,184),(92,160,87,184),(92,5,87,184),(210,5,87,184),(210,123,87,184),(210,13,87,184),(210,13,87,97),(210,13,87,104),(210,243,87,104),(210,243,128,104),(210,243,129,104),(5,243,129,104),(0,0,0,18),(0,0,125,18),(0,0,168,18),(0,0,221,18),(0,0,0,57),(167,0,0,57),(167,0,127,57),(217,0,127,57),(217,0,127,81),(217,0,127,208),(194,0,127,208),(194,0,199,208),(194,0,29,208),(130,0,29,208),(130,245,29,208),(10,245,29,208),(10,245,206,208),(10,245,146,208),(10,245,146,128),(165,245,146,128),(165,245,146,224),(165,245,146,33),(165,219,146,33),(165,219,146,212),(165,219,142,212),(165,219,142,128),(165,219,142,63),(165,161,142,63),(165,77,142,63),(165,185,142,63),(10,185,142,63),(142,185,142,63),(134,185,142,63),(0,0,104,0),(0,0,98,0),(6,0,98,0),(6,112,98,0),(6,55,98,0),(6,55,98,222),(6,234,98,222),(6,234,98,88),(6,203,98,88),(6,224,98,88),(120,224,98,88),(120,224,98,147),(120,9,98,147),(46,9,98,147),(46,9,166,147),(46,158,166,147),(46,158,166,250),(46,107,166,250),(46,107,108,250),(46,107,108,232),(46,107,123,232),(46,235,123,232),(46,57,123,232),(68,57,123,232),(68,57,123,115),(68,57,221,115),(68,57,71,115),(68,57,18,115),(68,57,18,187),(68,57,18,120),(0,0,206,0),(0,0,0,21),(33,0,0,21),(33,0,0,197),(123,0,0,197),(123,0,0,193),(123,0,0,4),(69,0,0,4),(69,0,0,229),(69,0,0,247),(69,0,101,247),(109,0,101,247),(109,0,101,112),(109,0,109,112),(109,7,109,112),(109,7,35,112),(109,7,35,209),(0,15,0,0),(0,0,74,0),(0,97,0,0),(147,97,0,0),(33,97,0,0),(33,83,0,0),(33,83,0,84),(33,83,136,84),(33,83,119,84),(33,36,119,84),(33,85,119,84),(33,85,126,84),(33,85,191,84),(33,85,191,20),(33,85,23,20),(33,85,141,20),(188,85,141,20),(76,85,141,20),(76,85,244,20),(76,85,244,104),(76,201,244,104),(195,201,244,104),(195,139,244,104),(0,0,215,0),(0,0,215,155),(0,0,4,155),(0,0,47,155),(0,255,47,155),(0,255,47,72),(0,255,87,72),(19,255,87,72),(93,0,0,0),(93,19,0,0),(93,19,0,64),(93,19,0,2),(93,19,0,72),(92,19,0,72),(92,19,212,72),(83,19,212,72),(225,19,212,72),(156,19,212,72),(156,254,212,72),(156,254,96,72),(156,34,96,72),(156,55,96,72),(156,237,96,72),(156,236,96,72),(26,236,96,72),(26,236,96,192),(26,236,96,215),(196,236,96,215),(196,236,96,71),(0,0,0,246),(78,0,0,246),(78,222,0,246),(78,222,0,189),(41,0,0,0),(41,0,0,106),(41,139,0,106),(41,139,157,106),(139,139,157,106),(139,169,157,106),(139,169,240,106),(139,169,240,231),(162,0,0,0),(162,38,0,0),(162,38,7,0),(162,38,46,0),(250,0,0,0),(250,112,0,0),(250,112,0,16),(48,112,0,16),(48,112,0,243),(48,112,0,135),(232,112,0,135),(232,112,5,135),(232,112,5,201),(232,112,80,201),(227,112,80,201),(227,112,80,222),(227,112,80,234),(51,112,80,234),(115,112,80,234),(151,112,80,234),(151,112,17,234),(151,167,17,234),(151,167,32,234),(158,167,32,234),(85,167,32,234),(85,226,32,234),(85,226,144,234),(85,226,138,234),(85,31,138,234),(85,31,73,234),(85,31,73,132),(85,31,73,124),(85,31,166,124),(85,31,17,124),(85,31,14,124),(15,31,14,124),(15,31,119,124),(15,31,107,124),(15,31,107,236),(15,188,107,236),(15,165,107,236),(15,165,107,215),(5,165,107,215),(41,165,107,215),(41,215,107,215),(41,215,107,19),(41,215,10,19),(41,215,10,225),(41,215,10,176),(15,215,10,176),(15,197,10,176),(15,197,158,176),(15,197,246,176),(15,197,246,46),(15,231,246,46),(15,231,246,207),(0,0,130,0),(156,0,130,0),(0,0,86,0),(50,0,86,0),(0,0,0,144),(0,0,0,93),(0,0,191,93),(0,66,191,93),(0,0,22,0),(0,160,22,0),(0,160,235,0),(0,160,235,22),(0,48,235,22),(0,187,235,22),(0,14,0,0),(228,14,0,0),(228,14,41,0),(228,112,41,0),(47,112,41,0),(47,112,6,0),(23,112,6,0),(114,112,6,0),(114,112,6,140),(114,59,6,140),(132,59,6,140),(132,72,6,140),(132,28,6,140),(171,28,6,140),(171,28,6,192),(171,28,6,193),(171,219,6,193),(171,219,194,193),(0,141,0,0),(0,0,223,0),(0,0,223,64),(240,0,223,64),(240,122,223,64),(240,154,223,64),(116,154,223,64),(116,172,223,64),(116,172,44,64),(116,172,98,64),(116,117,98,64),(44,117,98,64),(44,141,98,64),(44,141,98,155),(44,141,118,155),(44,141,103,155),(193,141,103,155),(193,141,105,155),(85,141,105,155),(89,141,105,155),(218,141,105,155),(218,226,105,155),(218,28,105,155),(218,191,105,155),(218,191,105,248),(202,0,0,0),(191,0,0,0),(0,177,0,0),(0,177,210,0),(232,177,210,0),(232,177,210,99),(232,9,210,99),(232,9,210,62),(232,9,210,151),(232,9,210,190),(96,0,0,0),(224,0,0,0),(224,18,0,0),(224,18,0,227),(224,18,0,127),(224,162,0,127),(224,162,71,127),(224,162,71,88),(224,162,81,88),(224,162,89,88),(224,162,114,88),(151,162,114,88),(151,162,114,131),(236,162,114,131),(236,51,114,131),(236,111,114,131),(236,111,114,29),(229,111,114,29),(0,0,0,129),(0,0,34,129),(0,0,66,129),(18,0,66,129),(233,0,66,129),(0,182,0,0),(90,182,0,0),(90,182,0,95),(219,182,0,95),(219,182,25,95),(219,182,25,209),(54,182,25,209),(54,82,25,209),(54,138,25,209),(205,138,25,209),(205,138,25,62),(205,8,25,62),(205,8,20,62),(115,8,20,62),(115,8,20,96),(115,158,20,96),(115,158,89,96),(115,158,89,35),(140,158,89,35),(140,238,89,35),(140,238,89,136),(122,238,89,136),(240,238,89,136),(240,238,177,136),(149,238,177,136),(149,41,177,136),(51,0,0,0),(67,0,0,0),(210,0,0,0),(210,0,238,0),(24,0,238,0),(24,171,238,0),(24,171,21,0),(24,171,21,121),(24,214,21,121),(75,214,21,121),(77,214,21,121),(200,214,21,121),(109,214,21,121),(109,236,21,121),(33,236,21,121),(88,236,21,121),(39,236,21,121),(39,236,21,226),(107,236,21,226),(107,8,21,226),(107,180,21,226),(38,180,21,226),(38,180,21,19),(254,180,21,19),(254,180,21,143),(254,180,21,134),(254,180,21,17),(254,180,21,215),(254,181,21,215),(254,181,107,215),(159,181,107,215),(159,111,107,215),(159,254,107,215),(159,254,161,215),(0,250,0,0),(0,250,174,0),(0,250,18,0),(0,250,18,126),(0,23,18,126),(0,23,8,126),(0,183,8,126),(0,183,150,126),(10,183,150,126),(10,208,150,126),(0,0,0,9),(179,0,0,9),(179,0,0,252),(179,239,0,252),(179,239,0,63),(179,239,0,27),(179,27,0,27),(120,27,0,27),(21,27,0,27),(21,27,182,27),(0,228,0,0),(0,228,0,110),(0,228,0,155),(0,228,0,169),(0,228,173,169),(18,228,173,169),(106,228,173,169),(70,228,173,169),(0,0,0,155),(89,0,0,155),(36,0,0,155),(36,198,0,155),(36,198,0,38),(222,198,0,38),(222,229,0,38),(222,123,0,38),(222,123,0,159),(222,123,37,159),(222,123,37,34),(222,123,125,34),(0,0,0,74),(0,0,170,74),(107,0,170,74),(107,0,170,22),(107,12,170,22),(0,0,172,0),(0,0,172,116),(0,0,172,160),(0,0,172,112),(0,30,172,112),(0,225,172,112),(0,38,172,112),(0,38,172,200),(0,38,172,63),(14,38,172,63),(14,11,172,63),(82,11,172,63),(82,215,172,63),(82,23,172,63),(144,23,172,63),(144,7,172,63),(144,7,172,139),(252,7,172,139),(252,175,172,139),(119,175,172,139),(119,175,24,139),(119,175,183,139),(119,40,183,139),(119,141,183,139),(119,141,183,61),(171,141,183,61),(171,141,183,245),(171,141,221,245),(69,141,221,245),(69,141,221,175),(69,97,221,175),(69,97,221,139),(69,97,188,139),(69,97,188,188),(158,97,188,188),(158,97,188,31),(158,113,188,31),(158,113,203,31),(243,113,203,31),(0,239,0,0),(0,133,0,0),(0,133,0,168),(0,47,0,168),(0,228,0,168),(0,228,0,164),(0,228,83,164),(0,0,11,0),(0,0,215,0),(0,0,73,0),(0,0,0,222),(0,0,47,222),(0,0,47,14),(0,0,47,159),(0,151,47,159),(0,179,47,159),(0,231,0,0),(0,156,0,0),(148,0,0,0),(148,50,0,0),(148,50,0,153),(148,50,118,153),(148,50,93,153),(148,103,93,153),(148,103,122,153),(148,103,122,25),(51,103,122,25),(51,72,122,25),(51,72,122,41),(51,72,122,107),(247,72,122,107),(247,72,147,107),(247,72,151,107),(247,72,151,106),(247,72,151,216),(247,72,151,148),(247,72,153,148),(247,73,153,148),(247,73,153,137),(247,122,153,137),(243,122,153,137),(0,0,47,0),(0,77,47,0),(0,77,47,79),(0,77,47,118),(0,77,47,205),(0,0,0,54),(0,0,0,243),(0,0,0,104),(204,0,0,104),(0,20,0,0),(68,20,0,0),(68,20,0,251),(68,20,213,251),(68,20,63,251),(68,136,63,251),(68,136,63,80),(68,136,199,80),(68,136,60,80),(68,136,195,80),(68,136,52,80),(68,136,52,91),(68,143,52,91),(0,0,223,0),(196,0,223,0),(200,0,223,0),(200,60,223,0),(215,60,223,0),(215,110,223,0),(215,110,135,0),(39,0,0,0),(39,184,0,0),(39,255,0,0),(39,255,0,127),(39,255,0,142),(39,255,0,229),(39,255,98,229),(0,0,0,111),(0,0,0,222),(0,199,0,222),(0,199,134,222),(0,199,134,116),(0,199,134,18),(0,199,134,140),(212,199,134,140),(212,95,134,140),(212,79,134,140),(212,79,134,140),(0,0,115,0),(0,0,115,196),(0,0,158,196),(227,0,158,196),(227,104,158,196),(229,104,158,196),(26,104,158,196),(0,75,0,0),(0,75,61,0),(0,75,220,0),(0,182,0,0),(178,182,0,0),(178,182,147,0),(125,182,147,0),(125,151,147,0),(0,0,0,113),(0,124,0,0),(0,124,0,167),(0,124,108,167),(0,124,108,225),(0,124,81,225),(0,184,81,225),(0,10,81,225),(0,10,243,225),(78,10,243,225),(78,226,243,225),(4,226,243,225),(4,226,243,5),(4,32,243,5),(192,32,243,5),(192,69,243,5),(192,69,243,197),(192,69,168,197),(192,69,180,197),(192,69,56,197),(192,69,166,197),(121,69,166,197),(121,229,166,197),(4,229,166,197),(4,229,200,197),(4,229,22,197),(4,229,22,80),(4,112,22,80),(4,112,22,187),(4,112,67,187),(12,112,67,187),(96,112,67,187),(96,236,67,187),(96,236,67,36),(96,216,67,36),(76,216,67,36),(76,216,112,36),(76,216,169,36),(58,216,169,36),(0,0,22,0),(0,0,22,169),(144,0,22,169),(16,0,22,169),(16,0,3,169),(16,0,215,169),(123,0,215,169),(123,92,215,169),(143,92,215,169),(143,20,215,169),(143,20,134,169),(143,20,134,200),(143,20,133,200),(136,20,133,200),(136,249,133,200),(136,62,133,200),(136,62,133,149),(136,228,133,149),(136,209,133,149),(136,209,133,37),(136,209,143,37),(64,209,143,37),(64,209,143,135),(64,73,143,135),(64,73,143,2),(64,73,72,2),(64,122,72,2),(64,122,87,2),(64,122,87,189),(64,122,134,189),(64,122,71,189),(64,122,229,189),(0,251,0,0),(0,251,0,0),(0,251,0,68),(0,29,0,68),(0,102,0,68),(0,185,0,68),(0,185,252,68),(0,185,40,68),(0,68,40,68),(0,139,0,0),(193,139,0,0),(234,139,0,0),(234,32,0,0),(0,0,0,166),(0,179,0,166),(0,179,0,237),(0,179,223,237),(0,179,124,237),(0,179,124,253),(57,179,124,253),(57,179,124,10),(57,179,66,10),(57,179,182,10),(57,179,182,241),(57,179,48,241),(57,82,48,241),(117,82,48,241),(50,82,48,241),(50,82,48,240),(50,82,48,159),(50,82,77,159),(50,82,5,159),(50,67,5,159),(53,67,5,159),(53,103,5,159),(114,103,5,159),(114,236,5,159),(168,236,5,159),(168,236,67,159),(194,236,67,159),(194,255,67,159),(194,255,107,159),(194,137,107,159),(148,137,107,159),(148,137,107,248),(148,137,92,248),(19,137,92,248),(19,137,35,248),(19,137,35,70),(19,137,254,70),(19,47,254,70),(0,0,37,0),(0,0,135,0),(165,0,135,0),(95,0,135,0),(95,22,135,0),(240,22,135,0),(73,22,135,0),(73,69,135,0),(73,140,135,0),(54,140,135,0),(54,140,135,253),(54,140,135,177),(195,140,135,177),(195,3,135,177),(195,3,49,177),(195,3,200,177),(195,3,220,177),(145,3,220,177),(145,3,220,230),(145,3,220,130),(145,3,27,130),(145,3,190,130),(0,0,35,0),(0,11,35,0),(0,11,35,209),(0,11,185,209),(78,11,185,209),(78,123,185,209),(207,123,185,209),(207,13,185,209),(207,13,185,48),(207,13,10,48),(207,13,255,48),(207,13,255,109),(207,61,255,109),(207,163,255,109),(207,31,255,109),(207,37,255,109),(207,37,66,109),(207,37,205,109),(207,214,205,109),(207,214,117,109),(207,214,129,109),(207,192,129,109),(207,192,63,109),(207,192,63,51),(207,193,63,51),(207,193,251,51),(29,193,251,51),(29,193,251,88),(29,193,211,88),(141,193,211,88),(141,193,112,88),(0,240,0,0),(186,240,0,0),(186,240,219,0),(186,240,219,173),(12,240,219,173),(12,198,219,173),(0,0,215,0),(0,0,215,201),(107,0,215,201),(255,0,215,201),(192,0,0,0),(192,0,0,251),(192,213,0,251),(192,213,228,251),(192,206,228,251),(0,0,132,0),(0,176,132,0),(0,176,132,98),(0,79,132,98),(0,79,132,231),(0,51,132,231),(0,51,222,231),(0,51,198,231),(0,0,198,231),(0,0,54,231),(127,0,54,231),(217,0,54,231),(217,0,155,231),(217,0,155,220),(217,33,155,220),(217,33,228,220),(217,33,81,220),(217,33,81,96),(0,0,246,0),(118,0,0,0),(118,0,164,0),(118,102,164,0),(118,102,56,0),(118,126,56,0),(118,126,120,0),(118,126,150,0),(118,126,109,0),(0,189,0,0),(0,189,0,93),(0,127,0,93),(0,127,0,250),(0,127,0,254),(0,127,0,38),(109,127,0,38),(105,127,0,38),(105,127,197,38),(105,191,197,38),(105,101,197,38),(105,172,197,38),(105,221,197,38),(197,221,197,38),(197,116,197,38),(197,116,197,215),(197,245,197,215),(139,245,197,215),(139,250,197,215),(25,250,197,215),(25,229,197,215),(25,229,197,222),(0,66,0,0),(0,66,45,0),(0,66,187,0),(0,177,187,0),(0,177,187,111),(0,177,228,111),(212,177,228,111),(227,177,228,111),(0,0,0,72),(0,0,0,70),(189,0,0,70),(78,0,0,70),(195,0,0,70),(195,199,0,70),(195,199,0,139),(119,199,0,139),(145,199,0,139),(176,199,0,139),(176,54,0,139),(176,245,0,139),(128,245,0,139),(0,0,0,167),(0,0,0,180),(0,0,241,180),(0,0,241,201),(0,0,51,201),(0,0,89,201),(0,0,89,181),(0,0,70,181),(0,179,70,181),(0,179,13,181),(0,64,13,181),(0,27,13,181),(0,27,13,82),(0,241,0,0),(172,241,0,0),(23,241,0,0),(23,176,0,0),(23,11,0,0),(23,11,0,219),(200,11,0,219),(200,11,0,250),(200,226,0,250),(200,226,46,250),(200,226,182,250),(200,82,182,250),(200,52,182,250),(126,52,182,250),(126,48,182,250),(0,0,206,0),(41,0,206,0),(41,0,244,0),(187,0,244,0),(187,0,244,0),(106,0,244,0),(106,0,244,179),(106,0,244,84),(57,0,244,84),(57,142,244,84),(57,227,244,84),(57,227,184,84),(54,227,184,84),(54,227,23,84),(167,227,23,84),(167,227,23,74),(167,227,23,154),(167,227,238,154),(167,227,238,193),(167,151,238,193),(167,119,238,193),(33,119,238,193),(33,119,238,177),(33,119,238,73),(33,217,238,73),(33,119,238,73),(33,236,238,73),(33,236,238,251),(160,236,238,251),(160,236,238,233),(160,236,238,160),(241,236,238,160),(241,236,238,252),(241,236,238,186),(241,236,238,177),(241,204,238,177),(241,174,238,177),(241,174,238,187),(241,174,238,193),(82,174,238,193),(247,174,238,193),(247,174,238,253),(247,174,238,186),(247,174,238,237),(247,174,252,237),(247,26,252,237),(247,182,252,237),(247,182,33,237),(135,182,33,237),(135,182,33,4),(135,182,33,73),(135,182,33,42),(13,182,33,42),(109,182,33,42),(115,182,33,42),(0,38,0,0),(12,38,0,0),(12,146,0,0),(12,131,0,0),(12,131,37,0),(12,43,37,0),(12,231,37,0),(12,231,37,215),(79,231,37,215),(79,213,37,215),(79,213,30,215),(79,213,15,215),(79,213,70,215),(0,0,0,57),(0,21,0,57),(0,21,0,230),(0,156,0,230),(0,123,0,230),(0,123,16,230),(0,123,16,242),(0,123,16,24),(0,123,16,13),(0,123,148,13),(0,123,37,13),(0,250,37,13),(0,250,56,13),(0,250,5,13),(166,250,5,13),(166,250,5,22),(166,250,5,170),(166,250,5,125),(0,0,0,117),(0,0,0,104),(1,0,0,104),(60,0,0,104),(60,0,0,179),(50,0,0,179),(50,0,66,179),(50,0,66,254),(50,0,118,254),(50,0,118,174),(141,0,118,174),(105,0,118,174),(105,55,118,174),(39,55,118,174),(92,55,118,174),(92,55,13,174),(149,55,13,174),(149,55,108,174),(149,244,108,174),(0,174,0,0),(0,174,0,176),(2,174,0,176),(2,233,0,176),(2,9,0,176),(2,9,0,130),(158,9,0,130),(158,9,0,0),(158,9,61,0),(158,9,126,0),(0,77,0,0),(0,0,0,72),(154,0,0,72),(154,0,0,54),(154,111,0,54),(154,111,0,25),(94,111,0,25),(94,134,0,25),(90,134,0,25),(90,230,0,25),(2,230,0,25),(77,230,0,25),(77,230,236,25),(77,230,236,49),(77,230,236,61),(128,230,236,61),(128,230,152,61),(39,230,152,61),(39,77,152,61),(39,77,179,61),(39,62,179,61),(87,62,179,61),(91,62,179,61),(91,62,179,78),(91,160,179,78),(91,160,179,48),(91,187,179,48),(187,187,179,48),(187,187,176,48),(0,57,0,0),(0,80,0,0),(254,80,0,0),(234,80,0,0),(136,0,0,0),(212,0,0,0),(212,0,0,96),(212,0,0,66),(212,0,0,184),(212,0,107,184),(247,0,107,184),(247,59,107,184),(247,237,107,184),(247,237,98,184),(195,237,98,184),(0,0,10,0),(0,28,10,0),(0,28,10,99),(0,30,10,99),(0,30,10,67),(0,158,10,67),(0,158,13,67),(0,158,27,67),(0,50,27,67),(0,50,27,129),(0,50,27,18),(0,249,27,18),(0,249,30,18),(0,249,30,245),(0,249,30,187),(166,249,30,187),(182,249,30,187),(182,249,30,38),(182,195,30,38),(182,195,30,243),(182,51,30,243),(182,51,65,243),(182,51,65,139),(182,51,128,139),(120,51,128,139),(232,51,128,139),(0,0,0,236),(0,192,0,236),(239,192,0,236),(0,221,0,0),(0,4,0,0),(0,4,159,0),(0,4,159,23),(52,4,159,23),(153,4,159,23),(153,239,159,23),(0,0,0,217),(0,203,0,217),(0,73,0,217),(0,191,0,217),(0,191,0,56),(137,0,0,0),(137,31,0,0),(137,31,146,0),(240,31,146,0),(240,31,62,0),(240,31,4,0),(113,31,4,0),(0,238,0,0),(191,238,0,0),(14,238,0,0),(211,238,0,0),(109,238,0,0),(109,177,0,0),(109,177,0,226),(109,177,190,226),(109,177,190,91),(109,190,190,91),(109,190,190,221),(109,190,197,221),(109,193,197,221),(109,193,197,202),(0,0,0,149),(102,0,0,149),(51,0,0,0),(100,0,0,0),(100,0,0,196),(100,0,0,69),(100,0,95,69),(237,0,0,0),(8,0,0,0),(8,0,0,202),(8,0,60,202),(0,0,40,0),(0,0,40,162),(0,188,0,0),(118,188,0,0),(118,170,0,0),(118,170,119,0),(0,83,0,0),(0,2,0,0),(0,2,208,0),(235,2,208,0),(202,2,208,0),(202,22,208,0),(188,22,208,0),(188,22,49,0),(131,22,49,0),(131,22,36,0),(206,22,36,0),(206,22,232,0),(171,22,232,0),(105,22,232,0),(105,22,184,0),(0,0,0,0),(172,0,0,0),(205,0,0,0),(78,0,0,0),(78,217,0,0),(78,127,0,0),(78,183,0,0),(78,52,0,0),(78,206,0,0),(78,206,0,194),(78,206,0,102),(78,85,0,102),(78,53,0,102),(78,82,0,102),(78,82,0,217),(78,82,0,237),(78,82,69,237),(78,20,69,237),(78,20,215,237),(78,20,215,191),(0,0,6,0),(0,0,0,229),(0,0,238,229),(0,0,238,78),(143,0,238,78),(107,0,238,78),(107,145,238,78),(174,145,238,78),(174,145,146,78),(249,145,146,78),(249,145,146,78),(249,145,108,78),(249,53,108,78),(249,53,108,203),(249,53,94,203),(249,53,200,203),(249,53,238,203),(249,53,178,203),(249,53,143,203),(249,53,180,203),(172,53,180,203),(172,139,180,203),(172,241,180,203),(172,242,180,203),(172,242,180,203),(246,242,180,203),(246,242,180,180),(246,242,180,188),(246,247,180,188),(72,247,180,188),(194,247,180,188),(194,247,180,45),(194,247,180,54),(30,0,0,0),(30,0,0,239),(30,0,3,239),(30,0,3,47),(30,0,152,47),(30,0,152,77),(30,0,189,77),(30,0,189,163),(30,0,189,159),(30,0,165,159),(89,0,0,0),(89,0,94,0),(89,0,94,0),(89,0,20,0),(140,0,0,0),(140,0,98,0),(140,0,212,0),(230,0,212,0),(230,0,105,0),(230,0,105,202),(0,146,0,0),(0,146,0,244),(0,227,0,0),(101,227,0,0),(101,227,0,32),(136,227,0,32),(136,227,148,32),(226,227,148,32),(226,227,148,17),(73,227,148,17),(162,227,148,17),(162,227,243,17),(162,227,93,17),(162,143,93,17),(162,143,93,246),(152,143,93,246),(152,143,177,246),(152,24,177,246),(54,24,177,246),(54,24,22,246),(54,24,22,108),(0,0,197,0),(0,0,197,100),(186,0,197,100),(50,0,197,100),(50,0,45,100),(50,231,45,100),(50,81,45,100),(30,81,45,100),(227,81,45,100),(227,81,96,100),(227,190,96,100),(227,190,96,54),(0,0,34,0),(0,0,235,0),(0,0,235,85),(0,105,235,85),(130,105,235,85),(130,16,235,85),(157,16,235,85),(157,16,242,85),(157,16,242,124),(157,253,242,124),(157,79,242,124),(157,126,242,124),(157,126,241,124),(157,126,167,124),(157,126,167,64),(157,126,167,120),(157,126,167,54),(157,65,167,54),(157,35,167,54),(157,35,101,54),(157,35,128,54),(157,148,128,54),(157,148,128,41),(157,189,128,41),(157,48,128,41),(0,0,0,1),(0,64,0,1),(0,64,0,23),(0,64,0,115),(0,139,0,115),(0,139,0,127),(71,139,0,127),(71,139,0,13),(166,139,0,13),(166,87,0,13),(166,87,0,214),(99,87,0,214),(99,87,79,214),(99,87,79,50),(99,170,79,50),(99,170,79,105),(99,170,79,105),(99,170,106,105),(99,170,106,92),(47,170,106,92),(64,170,106,92),(64,170,106,170),(111,170,106,170),(111,170,106,100),(111,170,131,100),(111,170,48,100),(237,0,0,0),(237,52,0,0),(0,0,126,0),(0,156,126,0),(0,200,126,0),(149,200,126,0),(149,83,126,0),(149,83,190,0),(149,83,190,102),(81,83,190,102),(50,83,190,102),(230,83,190,102),(230,219,190,102),(0,5,0,0),(0,5,91,0),(2,5,91,0),(2,5,60,0),(0,179,0,0),(0,179,0,170),(0,179,147,170),(142,0,0,0),(142,0,157,0),(146,0,157,0),(174,0,157,0),(174,92,157,0),(235,92,157,0),(235,92,157,191),(235,92,157,218),(235,92,157,116),(151,92,157,116),(151,88,157,116),(151,88,213,116),(151,88,207,116),(151,221,207,116),(151,221,168,116),(151,221,109,116),(151,221,109,222),(151,117,109,222),(151,132,109,222),(95,132,109,222),(95,132,40,222),(95,180,40,222),(95,37,40,222),(48,37,40,222),(179,37,40,222),(179,37,40,159),(179,37,147,159),(179,37,146,159),(4,37,146,159),(4,74,146,159),(4,74,3,159),(4,195,3,159),(4,195,12,159),(4,195,12,245),(4,195,12,227),(4,195,145,227),(4,197,145,227),(0,129,0,0),(184,129,0,0),(184,129,0,167),(82,129,0,167),(82,154,0,167),(82,125,0,167),(82,39,0,167),(82,39,22,167),(121,39,22,167),(121,39,216,167),(121,39,146,167),(74,39,146,167),(74,39,146,236),(0,224,0,0),(20,224,0,0),(191,224,0,0),(191,224,0,5),(191,224,231,5),(0,68,0,0),(117,68,0,0),(117,68,0,187),(117,68,0,105),(117,68,0,157),(80,68,0,157),(0,222,0,0),(0,219,0,0),(104,219,0,0),(104,219,195,0),(253,219,195,0),(253,219,148,0),(253,219,148,85),(253,82,148,85),(253,82,72,85),(0,247,0,0),(0,191,0,0),(0,238,0,0),(0,238,63,0),(0,230,63,0),(0,230,63,123),(0,230,63,135),(0,230,19,135),(23,230,19,135),(23,80,19,135),(23,80,19,150),(23,63,19,150),(23,63,213,150),(23,63,213,65),(23,63,211,65),(23,237,211,65),(23,237,211,78),(23,47,211,78),(23,47,8,78),(23,47,160,78),(23,47,160,70),(23,47,29,70),(23,47,29,81),(23,54,29,81),(23,54,112,81),(0,201,0,0),(174,201,0,0),(174,250,0,0),(174,250,60,0),(0,0,232,0),(0,0,128,0),(0,195,128,0),(0,113,128,0),(0,113,128,230),(0,100,128,230),(0,147,128,230),(0,222,128,230),(0,0,99,0),(224,0,99,0),(224,0,79,0),(224,0,208,0),(224,0,194,0),(94,0,194,0),(94,108,194,0),(98,0,0,0),(98,0,58,0),(98,0,32,0),(98,0,46,0),(98,184,46,0),(74,184,46,0),(74,184,46,110),(74,184,35,110),(74,116,35,110),(74,116,182,110),(74,188,182,110),(74,188,167,110),(74,2,167,110),(74,2,167,237),(36,2,167,237),(37,2,167,237),(156,2,167,237),(8,2,167,237),(8,2,170,237),(0,0,125,0),(0,0,125,239),(0,116,125,239),(0,116,125,40),(0,116,180,40),(129,116,180,40),(240,116,180,40),(216,116,180,40),(140,116,180,40),(0,10,0,0),(0,134,0,0),(0,134,39,0),(0,134,9,0),(0,104,9,0),(0,104,136,0),(0,104,107,0),(0,104,107,199),(0,104,188,199),(0,104,20,199),(0,25,20,199),(173,25,20,199),(173,19,20,199),(173,19,20,188),(173,19,20,86),(173,19,235,86),(173,19,235,84),(68,19,235,84),(54,19,235,84),(204,19,235,84),(204,19,192,84),(0,0,0,194),(0,0,0,194),(174,0,0,194),(174,0,253,194),(71,0,253,194),(71,15,253,194),(71,15,172,194),(200,0,0,0),(126,0,0,0),(126,254,0,0),(126,254,122,0),(126,112,122,0),(251,112,122,0),(182,112,122,0),(182,112,122,71),(182,112,122,112),(182,112,122,51),(182,92,122,51),(19,92,122,51),(19,92,122,3),(133,92,122,3),(199,92,122,3),(199,136,122,3),(111,136,122,3),(111,136,239,3),(111,136,239,3),(111,136,239,37),(111,136,239,80),(111,136,73,80),(111,136,73,109),(111,136,46,109),(156,136,46,109),(86,136,46,109),(163,0,0,0),(163,0,166,0),(61,0,166,0),(250,0,166,0),(40,0,166,0),(155,0,166,0),(212,0,0,0),(240,0,0,0),(240,0,147,0),(240,56,147,0),(0,0,0,110),(0,0,0,234),(0,0,0,106),(0,0,83,106),(18,0,0,0),(18,0,0,15),(18,0,0,239),(18,253,0,239),(18,253,177,239),(18,253,177,194),(0,0,68,0),(0,176,68,0),(105,176,68,0),(62,176,68,0),(100,176,68,0),(23,176,68,0),(23,176,22,0),(23,176,50,0),(23,254,50,0),(23,254,50,24),(23,254,52,24),(23,254,35,24),(51,254,35,24),(51,254,55,24),(125,254,55,24),(125,39,55,24),(37,39,55,24),(37,39,98,24),(37,217,98,24),(37,217,98,240),(37,8,98,240),(37,8,191,240),(37,101,191,240),(204,101,191,240),(204,55,191,240),(187,55,191,240),(187,55,191,123),(187,55,31,123),(187,114,31,123),(187,114,150,123),(187,114,150,59),(187,114,150,193),(187,114,150,38),(187,114,150,85),(187,114,14,85),(187,127,14,85),(0,0,156,0),(0,0,208,0),(0,0,208,225),(0,127,208,225),(0,127,208,46),(0,127,66,46),(0,168,66,46),(0,168,66,138),(227,168,66,138),(227,168,162,138),(99,168,162,138),(99,168,162,172),(99,10,162,172),(0,93,0,0),(46,93,0,0),(199,93,0,0),(199,93,198,0),(199,93,198,143),(199,93,247,143),(212,93,247,143),(57,93,247,143),(108,93,247,143),(108,82,247,143),(0,214,0,0),(197,214,0,0),(197,114,0,0),(197,149,0,0),(55,149,0,0),(55,149,0,106),(35,149,0,106),(35,149,0,158),(35,149,181,158),(35,59,181,158),(35,59,181,1),(35,118,181,1),(35,118,152,1),(35,118,152,75),(35,118,152,57),(35,118,208,57),(35,82,208,57),(35,82,208,57),(35,159,208,57),(35,159,233,57),(35,159,233,232),(35,159,193,232),(4,159,193,232),(107,159,193,232),(229,159,193,232),(229,159,193,200),(229,159,129,200),(204,159,129,200),(204,217,129,200),(204,217,73,200),(63,217,73,200),(63,217,73,102),(63,217,18,102),(63,217,18,31),(63,217,48,31),(0,0,0,226),(0,0,0,87),(80,0,0,87),(158,0,0,87),(158,6,0,87),(72,6,0,87),(72,6,0,101),(107,6,0,101),(107,6,41,101),(107,224,41,101),(107,150,41,101),(107,150,41,165),(107,95,41,165),(107,95,41,19),(107,95,41,46),(107,95,250,46),(0,0,0,38),(0,170,0,38),(0,170,0,67),(0,170,0,210),(0,170,0,82),(0,170,0,82),(0,0,0,176),(234,0,0,176),(234,150,0,176),(234,150,220,176),(0,97,0,0),(67,97,0,0),(67,241,0,0),(67,241,0,78),(67,26,0,78),(37,26,0,78),(40,0,0,0),(40,0,0,180),(204,0,0,180),(17,0,0,180),(17,181,0,180),(217,0,0,0),(0,0,0,220),(0,0,0,116),(0,0,0,18),(0,246,0,18),(0,28,0,18),(0,28,171,18),(0,28,171,24),(0,162,171,24),(202,162,171,24),(202,122,171,24),(202,122,152,24),(223,0,0,0),(223,233,0,0),(223,233,55,0),(48,233,55,0),(48,233,6,0),(0,0,0,171),(0,0,122,171),(0,0,122,214),(0,117,122,214),(0,11,122,214),(0,11,122,107),(0,11,31,107),(0,11,153,107),(0,11,214,107),(0,11,94,107),(0,11,57,107),(0,11,57,55),(0,11,57,24),(0,11,105,24),(0,11,82,24),(0,11,82,15),(0,244,82,15),(0,87,82,15),(0,121,82,15),(0,0,73,0),(0,205,73,0),(0,205,73,116),(0,205,119,116),(24,0,0,0),(105,0,0,0),(105,0,250,0),(88,0,250,0),(88,233,250,0),(88,233,43,0),(17,233,43,0),(17,185,43,0),(17,185,200,0),(17,19,200,0),(205,19,200,0),(40,19,200,0),(225,19,200,0),(138,0,0,0),(81,0,0,0),(81,0,0,151),(81,0,0,196),(105,0,0,196),(105,0,0,2),(1,0,0,2),(1,0,0,14),(1,0,0,170),(1,0,0,71),(1,0,60,71),(1,0,172,71),(34,0,172,71),(248,0,172,71),(134,0,172,71),(134,0,224,71),(134,0,224,179),(121,0,224,179),(121,160,224,179),(121,224,224,179),(0,17,0,0),(0,17,0,32),(238,17,0,32),(238,66,0,32),(238,218,0,32),(238,218,0,57),(238,116,0,57),(238,116,84,57),(238,116,185,57),(238,116,185,167),(238,139,185,167),(238,139,211,167),(238,139,183,167),(238,139,183,189),(238,139,59,189),(238,0,59,189),(238,0,59,240),(238,0,59,175),(238,0,54,175),(238,0,54,193),(238,0,54,24),(73,0,54,24),(73,138,54,24),(73,138,16,24),(73,138,193,24),(73,156,193,24),(0,0,0,185),(0,0,121,185),(159,0,121,185),(87,0,121,185),(0,195,0,0),(0,195,181,0),(0,195,175,0),(0,195,175,114),(0,99,175,114),(245,99,175,114),(124,99,175,114),(124,99,175,133),(124,99,22,133),(124,99,37,133),(124,118,37,133),(124,118,37,206),(124,118,216,206),(8,0,0,0),(102,0,0,0),(102,0,161,0),(102,0,161,131),(102,74,161,131),(102,74,161,244),(175,74,161,244),(175,74,161,87),(133,74,161,87),(182,74,161,87),(182,74,180,87),(182,74,180,120),(182,74,180,91),(182,74,244,91),(182,74,228,91),(211,74,228,91),(211,74,228,164),(211,213,228,164),(211,46,228,164),(211,46,228,141),(16,46,228,141),(16,83,228,141),(0,0,0,12),(211,0,0,12),(211,224,0,12),(211,224,44,12),(250,224,44,12),(17,224,44,12),(127,224,44,12),(127,224,153,12),(127,224,153,215),(127,61,153,215),(11,0,0,0),(11,10,0,0),(11,10,0,215),(74,10,0,215),(74,10,0,59),(74,10,0,15),(194,10,0,15),(194,10,102,15),(194,10,102,217),(194,10,102,1),(194,121,102,1),(194,121,102,44),(194,121,102,173),(194,121,102,15),(194,121,102,7),(194,8,102,7),(194,8,49,7),(194,8,49,95),(194,8,98,95),(194,11,98,95),(194,11,60,95),(194,166,60,95),(194,166,60,4),(194,166,175,4),(194,41,175,4),(194,41,173,4),(194,41,78,4),(194,41,78,97),(7,41,78,97),(7,41,22,97),(7,16,22,97),(7,16,22,115),(7,16,22,22),(0,0,246,0),(140,0,246,0),(140,0,246,123),(140,0,163,123),(140,203,163,123),(140,91,163,123),(140,91,163,24),(86,91,163,24),(86,152,163,24),(78,152,163,24),(78,19,163,24),(147,19,163,24),(147,63,163,24),(147,63,29,24),(147,216,29,24),(147,216,29,87),(147,216,9,87),(147,93,9,87),(147,93,171,87),(0,162,0,0),(49,162,0,0),(49,162,96,0),(128,162,96,0),(128,162,215,0),(128,162,124,0),(128,162,146,0),(128,68,146,0),(74,68,146,0),(74,106,146,0),(227,106,146,0),(227,38,146,0),(0,0,78,0),(0,0,246,0),(0,8,0,0),(0,8,119,0),(65,8,119,0),(57,8,119,0),(57,8,103,0),(57,118,103,0),(57,118,103,87),(138,0,0,0),(138,0,0,97),(138,0,0,236),(138,0,0,134),(186,0,0,134),(64,0,0,134),(64,0,0,137),(64,74,0,137),(64,173,0,137),(64,4,0,137),(64,4,0,140),(106,4,0,140),(61,4,0,140),(61,4,0,52),(187,4,0,52),(234,4,0,52),(234,4,0,123),(11,0,0,0),(11,80,0,0),(11,33,0,0),(0,107,0,0),(0,107,204,0),(29,107,204,0),(29,107,35,0),(29,107,90,0),(29,107,76,0),(29,107,174,0),(0,0,0,249),(0,0,9,249),(0,0,9,132),(0,0,135,132),(0,5,135,132),(0,5,135,210),(0,5,219,210),(0,5,219,109),(0,69,0,0),(168,69,0,0),(168,69,171,0),(168,69,171,240),(30,69,171,240),(30,208,171,240),(30,205,171,240),(30,205,24,240),(30,205,240,240),(210,0,0,0),(210,110,0,0),(210,110,0,250),(51,110,0,250),(51,110,51,250),(51,110,51,232),(51,110,51,144),(64,110,51,144),(64,110,51,164),(209,110,51,164),(209,110,51,138),(209,110,246,138),(209,110,131,138),(209,106,131,138),(130,106,131,138),(130,106,225,138),(130,253,225,138),(130,253,172,138),(130,253,28,138),(130,253,96,138),(130,223,96,138),(130,252,96,138),(91,252,96,138),(91,222,96,138),(0,36,0,0),(5,36,0,0),(5,36,0,160),(5,60,0,160),(5,60,0,254),(5,60,0,93),(5,60,0,126),(5,60,0,225),(5,29,0,225),(5,75,0,225),(101,75,0,225),(251,75,0,225),(251,248,0,225),(148,248,0,225),(148,155,0,225),(148,71,0,225),(148,232,0,225),(148,246,0,225),(51,246,0,225),(51,246,225,225),(51,246,104,225),(0,161,0,0),(0,161,222,0),(0,161,59,0),(0,161,127,0),(220,161,127,0),(220,16,127,0),(220,16,127,46),(220,16,127,48),(58,16,127,48),(58,232,127,48),(0,0,0,175),(100,0,0,175),(100,216,0,175),(167,216,0,175),(144,216,0,175),(144,216,12,175),(58,216,12,175),(39,216,12,175),(12,216,12,175),(107,216,12,175),(107,216,12,62),(107,216,12,2),(107,216,12,38),(107,195,12,38),(107,195,231,38),(107,38,231,38),(107,170,231,38),(107,170,231,35),(107,223,231,35),(107,223,236,35),(107,223,246,35),(255,223,246,35),(0,0,0,0),(0,0,0,235),(0,20,0,235),(70,20,0,235),(70,133,0,235),(70,133,0,66),(70,133,0,137),(219,0,0,0),(178,0,0,0),(178,0,174,0),(44,0,174,0),(0,194,0,0),(0,194,116,0),(0,194,116,98),(219,194,116,98),(219,194,116,104),(219,194,116,82),(236,194,116,82),(76,0,0,0),(57,0,0,0),(0,0,209,0),(0,0,209,30),(0,0,209,235),(0,0,192,235),(0,0,192,253),(0,138,192,253),(177,138,192,253),(177,138,192,207),(177,138,40,207),(177,138,40,158),(107,0,0,0),(159,0,0,0),(0,0,0,53),(0,210,0,53),(0,210,29,53),(0,5,29,53),(0,5,29,85),(0,30,29,85),(0,30,67,85),(0,238,67,85),(0,102,0,0),(0,133,0,0),(0,133,0,163),(0,22,0,163),(118,22,0,163),(118,22,0,27),(118,22,205,27),(118,22,100,27),(118,22,56,27),(118,22,56,82),(45,22,56,82),(108,22,56,82),(108,22,14,82),(108,140,14,82),(108,140,14,249),(108,86,14,249),(108,133,14,249),(108,133,14,17),(124,133,14,17),(120,133,14,17),(44,133,14,17),(44,133,14,219),(44,133,14,140),(44,178,14,140),(44,178,14,67),(44,134,14,67),(44,101,14,67),(44,101,89,67),(44,101,192,67),(44,101,56,67),(66,101,56,67),(66,101,70,67),(66,101,70,99),(66,101,106,99),(141,101,106,99),(141,101,106,15),(65,0,0,0),(63,0,0,0),(63,207,0,0),(63,207,17,0),(63,207,209,0),(36,0,0,0),(36,67,0,0),(195,67,0,0),(195,237,0,0),(0,229,0,0),(180,229,0,0),(0,97,0,0),(0,0,85,0),(0,61,85,0),(0,127,85,0),(190,127,85,0),(3,127,85,0),(3,127,207,0),(3,127,64,0),(3,104,64,0),(3,104,64,235),(3,104,64,250),(3,104,18,250),(0,13,0,0),(0,13,146,0),(0,13,146,178),(160,13,146,178),(124,13,146,178),(124,77,146,178),(225,77,146,178),(225,24,146,178),(225,204,146,178),(121,204,146,178),(121,204,146,58),(121,204,229,58),(121,204,101,58),(10,204,101,58),(0,0,0,68),(0,124,0,68),(0,253,0,68),(0,253,0,124),(255,0,0,0),(112,0,0,0),(112,244,0,0),(112,244,0,80),(198,244,0,80),(198,126,0,80),(198,126,8,80),(198,127,8,80),(198,127,8,215),(0,19,0,0),(0,19,78,0),(21,0,0,0),(21,0,0,18),(21,0,136,18),(21,36,136,18),(21,36,136,75),(21,36,136,198),(21,36,136,171),(21,125,136,171),(21,125,148,171),(21,125,148,7),(245,125,148,7),(245,213,148,7),(198,213,148,7),(4,213,148,7),(4,118,148,7),(4,88,148,7),(4,88,216,7),(252,88,216,7),(252,175,216,7),(252,117,216,7),(0,171,0,0),(0,171,99,0),(0,171,25,0),(0,171,25,104),(0,171,25,198),(0,63,25,198),(0,63,93,198),(146,63,93,198),(146,63,93,221),(146,63,93,196),(146,63,93,190),(146,12,93,190),(146,86,93,190),(146,86,93,94),(0,160,0,0),(0,160,10,0),(0,160,10,102),(213,160,10,102),(213,160,251,102),(0,152,0,0),(0,152,0,105),(0,110,0,105),(252,110,0,105),(252,110,0,66),(218,0,0,0),(0,0,0,0),(0,0,0,195),(0,0,0,230),(249,0,0,230),(249,0,0,99),(249,21,0,99),(38,21,0,99),(38,120,0,99),(48,120,0,99),(48,120,200,99),(11,120,200,99),(11,120,170,99),(79,0,0,0),(79,157,0,0),(79,247,0,0),(151,247,0,0),(151,11,0,0),(86,0,0,0),(86,0,0,78),(86,0,92,78),(86,39,92,78),(86,221,92,78),(86,47,92,78),(86,156,92,78),(86,237,92,78),(86,237,92,165),(86,237,92,221),(86,74,92,221),(57,74,92,221),(57,136,92,221),(225,136,92,221),(197,136,92,221),(197,136,92,112),(169,136,92,112),(169,136,92,17),(0,0,0,90),(117,0,0,90),(117,0,0,114),(141,0,0,114),(226,0,0,114),(9,0,0,114),(9,0,224,114),(184,0,224,114),(184,0,14,114),(112,0,14,114),(112,0,112,114),(112,227,112,114),(112,197,112,114),(13,197,112,114),(13,197,141,114),(13,197,141,114),(166,197,141,114),(166,234,141,114),(166,234,241,114),(166,234,241,73),(166,234,195,73),(166,49,195,73),(166,197,195,73),(166,96,195,73),(166,43,195,73),(183,43,195,73),(64,43,195,73),(64,5,195,73),(64,5,195,192),(3,5,195,192),(3,241,195,192),(3,199,195,192),(0,48,0,0),(0,247,0,0),(0,0,173,0),(0,131,173,0),(172,131,173,0),(172,131,173,38),(172,71,173,38),(49,71,173,38),(204,71,173,38),(174,71,173,38),(174,73,173,38),(174,65,173,38),(142,65,173,38),(142,154,173,38),(142,154,155,38),(142,154,214,38),(142,154,214,118),(142,154,115,118),(142,73,115,118),(112,73,115,118),(0,0,187,0),(0,0,218,0),(0,14,218,0),(0,14,218,80),(0,14,243,80),(0,205,243,80),(0,205,52,80),(0,15,52,80),(0,15,27,80),(91,15,27,80),(91,15,112,80),(91,15,112,238),(0,0,0,18),(0,0,0,17),(0,233,0,17),(0,233,0,104),(0,52,0,104),(0,52,1,104),(205,52,1,104),(205,52,218,104),(205,52,218,235),(205,188,218,235),(205,245,218,235),(124,245,218,235),(124,245,218,121),(124,245,218,152),(124,123,218,152),(124,123,36,152),(124,123,36,236),(52,123,36,236),(52,123,100,236),(52,123,100,190),(52,14,100,190),(52,185,100,190),(52,185,128,190),(52,185,128,109),(52,185,128,236),(52,62,128,236),(52,26,128,236),(52,117,128,236),(52,117,128,98),(52,117,222,98),(52,117,89,98),(21,117,89,98),(138,117,89,98),(0,81,0,0),(0,81,4,0),(0,81,232,0),(0,81,232,248),(0,81,232,172),(0,81,82,172),(0,81,82,28),(154,81,82,28),(154,81,82,124),(161,0,0,0),(161,0,0,208),(0,0,1,0),(5,0,1,0),(5,0,10,0),(208,0,10,0),(142,0,10,0),(142,0,10,145),(142,221,10,145),(142,221,10,196),(142,26,10,196),(142,26,209,196),(142,26,52,196),(142,26,52,182),(142,26,52,183),(142,26,52,254),(142,26,52,100),(142,26,1,100),(0,63,0,0),(0,143,0,0),(0,143,247,0),(0,143,107,0),(191,143,107,0),(191,143,142,0),(191,143,142,247),(191,130,142,247),(223,130,142,247),(0,108,0,0),(242,108,0,0),(242,108,0,178),(242,238,0,178),(242,151,0,178),(0,0,104,0),(113,0,104,0),(113,0,104,7),(0,0,118,0),(0,0,118,149),(0,0,42,149),(125,0,42,149),(125,0,42,78),(125,0,42,152),(125,98,42,152),(125,98,42,143),(125,30,42,143),(125,30,42,254),(125,30,42,51),(125,167,42,51),(177,167,42,51),(177,167,117,51),(0,0,0,104),(188,0,0,104),(188,0,0,28),(95,0,0,28),(95,185,0,28),(109,185,0,28),(0,66,0,0),(0,58,0,0),(0,241,0,0),(138,241,0,0),(138,241,147,0),(138,241,147,79),(145,241,147,79),(145,241,24,79),(113,241,24,79),(0,0,8,0),(119,0,8,0),(119,0,199,0),(119,105,199,0),(0,152,0,0),(0,169,0,0),(95,0,0,0),(95,189,0,0),(95,189,125,0),(95,217,125,0),(0,0,0,216),(0,0,0,178),(0,0,78,178),(0,0,45,178),(0,62,45,178),(0,103,45,178),(0,83,45,178),(0,90,45,178),(0,52,45,178),(0,52,194,178),(0,21,194,178),(0,21,10,178),(0,21,190,178),(0,21,19,178),(0,168,19,178),(226,168,19,178),(228,168,19,178),(228,30,19,178),(104,30,19,178),(104,30,19,94),(218,30,19,94),(218,30,19,176),(218,30,19,120),(218,184,19,120),(218,184,1,120),(218,184,1,99),(218,184,51,99),(218,184,66,99),(218,13,66,99),(218,132,66,99),(218,132,39,99),(218,132,248,99),(218,132,58,99),(218,132,58,241),(218,132,58,239),(218,132,1,239),(218,132,158,239),(218,132,69,239),(218,132,107,239),(218,132,88,239),(176,132,88,239),(176,132,99,239),(176,23,99,239),(242,23,99,239),(116,23,99,239),(82,23,99,239),(141,23,99,239),(141,10,99,239),(73,10,99,239),(73,67,99,239),(43,67,99,239),(171,67,99,239),(171,67,45,239),(171,18,45,239),(171,96,45,239),(17,96,45,239),(17,173,45,239),(17,173,233,239),(88,173,233,239),(158,173,233,239),(0,0,0,143),(12,0,0,143),(217,0,0,143),(217,196,0,143),(217,5,0,143),(217,5,0,92),(217,5,176,92),(217,5,176,20),(217,5,176,174),(217,5,126,174),(38,5,126,174),(38,5,126,16),(136,5,126,16),(136,3,126,16),(136,3,150,16),(98,3,150,16),(98,3,7,16),(98,3,7,56),(98,3,7,93),(98,3,7,47),(51,0,0,0),(51,0,0,215),(51,0,0,115),(235,0,0,115),(216,0,0,115),(216,0,0,119),(235,0,0,119),(69,0,0,119),(69,0,31,119),(69,0,109,119),(69,89,109,119),(69,89,67,119),(69,144,67,119),(69,144,103,119),(69,144,86,119),(69,241,86,119),(69,29,86,119),(69,131,86,119),(144,131,86,119),(144,131,100,119),(214,131,100,119),(53,0,0,0),(214,0,0,0),(214,98,0,0),(214,40,0,0),(214,248,0,0),(214,248,125,0),(238,0,0,0),(238,0,122,0),(238,0,30,0),(238,0,62,0),(238,0,150,0),(238,191,150,0),(42,191,150,0),(226,191,150,0),(231,191,150,0),(204,191,150,0),(163,191,150,0),(118,191,150,0),(159,191,150,0),(159,191,39,0),(159,191,221,0),(167,191,221,0),(167,191,221,221),(167,29,221,221),(167,121,221,221),(167,178,221,221),(167,50,221,221),(167,50,67,221),(0,0,0,161),(0,0,0,35),(0,208,0,35),(68,208,0,35),(68,208,0,101),(0,253,0,0),(0,253,185,0),(0,0,0,85),(0,0,0,11),(0,0,0,152),(251,0,0,0),(251,0,202,0),(251,114,202,0),(251,168,202,0),(251,168,202,130),(251,7,202,130),(251,7,209,130),(41,7,209,130),(41,7,148,130),(41,7,148,137),(245,7,148,137),(245,7,203,137),(245,7,203,142),(245,113,203,142),(245,113,47,142),(245,113,47,190),(245,113,235,190),(245,113,139,190),(245,243,139,190),(59,243,139,190),(59,155,139,190),(126,155,139,190),(126,105,139,190),(126,187,139,190),(126,145,139,190),(126,179,139,190),(126,179,139,95),(126,218,139,95),(197,218,139,95),(197,218,139,153),(197,218,113,153),(197,112,113,153),(197,112,113,88),(79,112,113,88),(79,112,113,31),(79,112,187,31),(79,112,187,234),(79,112,187,42),(79,112,187,61),(36,0,0,0),(0,0,0,84),(0,196,0,84),(161,196,0,84),(161,196,13,84),(161,196,22,84),(161,196,248,84),(161,196,248,77),(161,196,253,77),(118,196,253,77),(118,196,253,26),(118,196,253,60),(0,0,0,160),(0,188,0,0),(0,188,0,0),(4,188,0,0),(4,167,0,0),(4,167,0,188),(4,167,0,34),(4,167,81,34),(4,167,81,230),(4,167,81,230),(95,167,81,230),(95,207,81,230),(95,159,81,230),(95,159,139,230),(95,159,139,164),(95,159,139,184),(95,175,139,184),(230,0,0,0),(167,0,0,0),(167,0,0,135),(0,0,90,0),(0,0,90,126),(0,202,90,126),(0,34,90,126),(0,34,104,126),(0,34,104,116),(0,34,222,116),(0,52,222,116),(0,52,188,116),(0,52,61,116),(0,57,61,116),(0,57,11,116),(25,57,11,116),(25,57,17,116),(69,57,17,116),(69,172,17,116),(69,120,17,116),(18,120,17,116),(50,120,17,116),(50,144,17,116),(0,0,222,0),(0,0,222,142),(0,0,222,115),(0,155,0,0),(0,155,226,0),(0,155,109,0),(0,224,109,0),(0,52,109,0),(0,52,109,201),(161,52,109,201),(161,150,109,201),(161,150,29,201),(0,64,0,0),(201,64,0,0),(201,153,0,0),(201,153,25,0),(0,0,24,0),(0,0,84,0),(0,0,45,0),(0,0,63,0),(84,0,63,0),(84,0,92,0),(84,0,97,0),(181,0,97,0),(181,0,97,85),(181,83,97,85),(4,0,0,0),(4,0,141,0),(0,0,63,0),(0,0,63,53),(240,0,63,53),(240,0,145,53),(152,0,145,53),(152,8,145,53),(152,212,145,53),(152,53,145,53),(152,53,28,53),(152,53,28,177),(152,95,28,177),(152,97,28,177),(69,97,28,177),(131,97,28,177),(107,97,28,177),(201,97,28,177),(201,163,28,177),(201,163,114,177),(201,163,114,43),(0,135,0,0),(241,135,0,0),(201,0,0,0),(201,0,150,0),(19,0,150,0),(19,0,197,0),(19,0,200,0),(19,0,200,240),(233,0,200,240),(233,0,200,156),(233,0,200,211),(233,197,200,211),(233,62,200,211),(0,0,0,164),(0,0,0,42),(49,0,0,42),(49,52,0,42),(49,253,0,42),(49,120,0,42),(49,120,0,221),(0,0,222,0),(0,58,222,0),(0,58,113,0),(0,58,113,81),(0,58,212,81),(0,149,212,81),(0,149,85,81),(0,149,92,81),(0,149,92,205),(87,149,92,205),(87,149,92,148),(87,149,92,4),(87,149,92,240),(87,149,211,240),(87,75,211,240),(13,75,211,240),(195,75,211,240),(64,75,211,240),(64,75,19,240),(4,0,0,0),(0,0,0,207),(49,0,0,207),(49,0,0,39),(0,184,0,0),(0,184,255,0),(0,160,255,0),(0,60,0,0),(0,60,0,161),(0,60,132,161),(0,154,132,161),(53,154,132,161),(0,0,96,0),(0,202,0,0),(0,202,165,0),(0,202,165,77),(0,202,165,248),(0,202,165,106),(0,202,165,154),(0,202,38,154),(0,71,38,154),(235,71,38,154),(235,71,83,154),(235,71,83,4),(235,160,83,4),(230,160,83,4),(230,160,178,4),(230,160,202,4),(230,160,131,4),(230,160,75,4),(230,160,206,4),(230,160,130,4),(0,0,0,201),(0,124,0,201),(0,124,0,85),(8,124,0,85),(8,127,0,85),(8,166,0,85),(8,155,0,85),(8,173,0,85),(8,80,0,85),(8,80,0,38),(8,80,0,42),(8,60,0,42),(8,173,0,42),(8,173,0,149),(8,173,138,149),(8,173,60,149),(8,173,60,131),(8,173,126,131),(8,173,154,131),(8,173,125,131),(19,173,125,131),(240,173,125,131),(0,0,20,0),(235,0,20,0),(235,0,112,0),(235,0,165,0),(235,0,106,0),(235,120,106,0),(235,120,106,121),(235,177,106,121),(235,177,242,121),(235,177,242,38),(235,177,215,38),(235,60,215,38),(235,60,215,222),(235,60,215,197),(0,0,78,0),(0,142,78,0),(0,28,78,0),(198,28,78,0),(198,163,78,0),(198,163,116,0),(241,163,116,0),(31,163,116,0),(31,163,116,67),(31,231,116,67),(31,227,116,67),(31,177,116,67),(31,8,116,67),(31,162,116,67),(31,162,116,212),(31,162,15,212),(4,162,15,212),(4,162,148,212),(140,162,148,212),(140,96,148,212),(140,96,148,99),(216,96,148,99),(0,0,0,10),(0,0,0,5),(0,93,0,5),(0,93,17,5),(0,93,17,89),(0,93,17,157),(162,93,17,157),(162,128,17,157),(162,128,230,157),(162,36,230,157),(183,36,230,157),(183,36,230,165),(176,36,230,165),(208,36,230,165),(208,36,55,165),(75,36,55,165),(38,36,55,165),(96,0,0,0),(96,225,0,0),(96,225,251,0),(96,148,251,0),(163,0,0,0),(163,181,0,0),(163,181,0,78),(163,181,0,173),(163,187,0,173),(0,188,0,0),(0,250,0,0),(0,250,0,194),(0,250,164,194),(0,171,164,194),(0,171,99,194),(0,235,99,194),(0,235,41,194),(14,235,41,194),(14,235,71,194),(14,235,71,57),(0,0,144,0),(0,0,94,0),(70,0,94,0),(70,0,94,154),(70,46,94,154),(70,46,94,139),(70,50,94,139),(93,50,94,139),(93,177,94,139),(93,177,94,198),(93,138,94,198),(93,116,94,198),(188,116,94,198),(188,123,94,198),(0,95,0,0),(0,144,0,0),(0,144,0,226),(0,144,0,113),(0,144,0,64),(0,144,152,64),(0,141,152,64),(0,205,0,0),(18,205,0,0),(50,205,0,0),(246,205,0,0),(246,205,0,189),(246,190,0,189),(246,190,77,189),(59,190,77,189),(59,200,77,189),(0,240,0,0),(73,240,0,0),(73,240,130,0),(73,240,11,0),(73,37,11,0),(73,37,11,132),(73,37,25,132),(22,37,25,132),(22,159,25,132),(31,159,25,132),(31,159,69,132),(31,133,69,132),(31,208,69,132),(116,208,69,132),(116,208,69,152),(52,208,69,152),(52,208,9,152),(52,194,9,152),(52,194,9,107),(52,194,9,228),(52,194,253,228),(52,194,135,228),(52,194,135,2),(52,194,63,2),(52,241,63,2),(52,241,63,120),(52,111,63,120),(52,161,63,120),(52,173,63,120),(52,173,39,120),(52,173,39,128),(52,173,169,128),(108,0,0,0),(108,0,0,213),(86,0,0,213),(223,0,0,213),(223,0,251,213),(223,239,251,213),(223,110,251,213),(223,110,251,115),(223,241,251,115),(223,241,130,115),(223,30,130,115),(0,0,0,188),(0,112,0,188),(0,112,0,86),(81,0,0,0),(81,12,0,0),(81,12,159,0),(81,12,159,209),(81,12,186,209),(81,12,169,209),(36,12,169,209),(142,0,0,0),(142,0,147,0),(142,0,147,184),(142,251,147,184),(241,251,147,184),(241,229,147,184),(241,229,147,101),(241,45,147,101),(241,45,147,9),(79,45,147,9),(79,45,147,165),(66,0,0,0),(66,252,0,0),(178,252,0,0),(178,15,0,0),(178,151,0,0),(178,151,179,0),(178,151,179,152),(122,0,0,0),(122,0,0,87),(122,0,0,166),(11,0,0,166),(11,0,0,188),(11,222,0,188),(11,222,0,105),(11,244,0,105),(137,0,0,0),(254,0,0,0),(0,0,223,0),(0,160,223,0),(0,0,0,97),(0,0,10,97),(0,0,10,146),(0,0,10,74),(54,0,10,74),(54,0,184,74),(112,0,184,74),(112,0,71,74),(112,0,246,74),(112,0,155,74),(3,0,155,74),(3,51,155,74),(3,51,8,74),(3,51,34,74),(3,87,34,74),(3,87,34,188),(3,87,22,188),(3,87,173,188),(3,87,4,188),(23,87,4,188),(23,87,200,188),(23,16,200,188),(23,57,200,188),(23,57,237,188),(23,156,237,188),(110,156,237,188),(110,166,237,188),(110,65,237,188),(0,16,0,0),(0,54,0,0),(0,50,0,0),(0,128,0,0),(0,177,0,0),(100,177,0,0),(100,59,0,0),(0,0,0,216),(26,0,0,216),(26,213,0,216),(26,213,0,33),(227,0,0,0),(227,194,0,0),(227,115,0,0),(227,33,0,0),(227,186,0,0),(227,186,0,3),(180,186,0,3),(180,186,145,3),(119,186,145,3),(119,186,145,115),(119,186,145,54),(119,186,145,221),(119,186,57,221),(119,158,57,221),(0,0,224,0),(0,79,224,0),(0,183,224,0),(203,183,224,0),(203,172,224,0),(203,172,58,0),(203,172,58,16),(203,170,58,16),(203,170,0,16),(203,170,166,16),(0,0,227,0),(104,0,227,0),(104,0,127,0),(104,24,127,0),(104,5,127,0),(104,5,159,0),(104,5,209,0),(57,5,209,0),(164,5,209,0),(164,5,209,89),(164,125,209,89),(164,125,118,89),(164,125,195,89),(167,125,195,89),(0,0,0,145),(0,0,0,50),(0,0,157,50),(0,44,157,50),(0,25,157,50),(10,25,157,50),(10,25,157,59),(10,25,157,27),(10,25,157,226),(10,25,41,226),(10,25,111,226),(10,25,89,226),(0,0,136,0),(0,91,136,0),(238,91,136,0),(238,91,136,122),(0,56,0,0),(164,56,0,0),(164,56,0,180),(164,200,0,180),(164,103,0,180),(164,151,0,180),(189,151,0,180),(189,151,213,180),(189,151,213,1),(189,151,213,156),(189,151,128,156),(65,151,128,156),(189,151,128,156),(130,151,128,156),(147,0,0,0),(147,0,0,20),(17,0,0,20),(17,115,0,20),(17,115,232,20),(17,115,100,20),(172,0,0,0),(172,0,0,97),(177,0,0,97),(177,0,186,97),(68,0,186,97),(68,0,155,97),(46,0,155,97),(46,150,155,97),(0,0,0,194),(0,16,0,194),(44,16,0,194),(44,162,0,194),(44,10,0,194),(44,10,201,194),(240,10,201,194),(0,0,0,8),(84,0,0,8),(84,0,0,183),(84,0,0,59),(84,0,183,59),(143,0,0,0),(143,0,0,125),(0,0,117,0),(147,0,117,0),(147,0,117,0),(147,0,117,211),(147,0,117,249),(0,11,0,0),(80,11,0,0),(80,11,125,0),(80,11,51,0),(80,11,51,217),(80,11,51,109),(197,11,51,109),(86,11,51,109),(86,11,4,109),(86,11,88,109),(86,249,88,109),(86,112,88,109),(86,112,88,54),(86,112,25,54),(86,112,116,54),(86,215,116,54),(86,215,180,54),(86,245,180,54),(53,245,180,54),(53,229,180,54),(53,102,180,54),(53,102,139,54),(53,102,139,132),(10,102,139,132),(10,102,118,132),(10,34,118,132),(10,34,157,132),(10,34,197,132),(10,34,139,132),(10,34,125,132),(21,0,0,0),(21,54,0,0),(21,214,0,0),(21,214,0,68),(21,253,0,68),(21,253,23,68),(21,253,23,0),(21,47,23,0),(21,47,23,72),(21,47,100,72),(206,47,100,72),(0,79,0,0),(19,79,0,0),(0,0,71,0),(0,0,71,239),(0,5,71,239),(0,5,11,239),(0,5,11,135),(224,5,11,135),(224,5,119,135),(224,5,119,154),(224,5,166,154),(224,5,166,255),(224,171,166,255),(224,171,166,134),(224,17,166,134),(18,0,0,0),(18,131,0,0),(18,131,195,0),(178,131,195,0),(178,131,206,0),(231,131,206,0),(231,57,206,0),(138,57,206,0),(254,57,206,0),(254,230,206,0),(20,230,206,0),(20,230,206,17),(20,230,206,205),(0,64,0,0),(0,64,0,85),(0,53,0,85),(0,53,0,194),(0,80,0,0),(0,80,193,0),(0,80,75,0),(81,80,75,0),(81,80,196,0),(81,80,220,0),(0,0,240,0),(0,0,26,0),(0,0,26,154),(218,0,26,154),(100,0,26,154),(100,21,26,154),(100,21,26,141),(0,80,0,0),(204,80,0,0),(204,80,0,17),(204,88,0,17),(204,87,0,17),(204,87,138,17),(204,87,138,191),(8,87,138,191),(8,20,138,191),(0,0,140,0),(124,0,140,0),(22,0,140,0),(22,212,140,0),(22,212,140,242),(22,212,140,115),(140,212,140,115),(111,212,140,115),(111,212,140,72),(111,129,140,72),(84,129,140,72),(84,129,169,72),(84,236,169,72),(151,236,169,72),(151,177,169,72),(151,63,169,72),(151,63,98,72),(151,63,98,97),(151,63,42,97),(151,63,199,97),(151,63,213,97),(151,63,145,97),(0,0,238,0),(0,0,250,0),(165,0,250,0),(165,0,250,135),(146,0,250,135),(146,0,250,184),(146,0,250,252),(34,0,250,252),(78,0,250,252),(164,0,250,252),(164,0,239,252),(164,75,239,252),(164,75,239,196),(164,75,208,196),(164,55,208,196),(164,55,79,196),(164,55,79,53),(164,55,151,53),(164,55,203,53),(164,25,203,53),(164,25,237,53),(164,25,182,53),(164,25,182,53),(193,25,182,53),(193,25,155,53),(199,25,155,53),(199,155,155,53),(132,155,155,53),(132,155,155,252),(132,36,155,252),(132,237,155,252),(132,237,155,29),(132,237,225,29),(132,237,225,53),(0,0,53,0),(0,0,159,0),(176,0,159,0),(0,180,0,0),(0,180,201,0),(0,180,192,0),(0,77,192,0),(0,77,30,0),(253,77,30,0),(223,77,30,0),(223,77,30,247),(223,77,30,130),(223,77,223,130),(223,77,69,130),(223,77,69,245),(123,77,69,245),(0,0,0,244),(0,0,175,244),(0,0,175,247),(0,0,210,247),(147,0,210,247),(147,0,210,174),(105,0,210,174),(105,0,210,131),(105,0,97,131),(105,22,97,131),(105,22,249,131),(254,22,249,131),(254,22,249,190),(254,22,14,190),(0,0,170,0),(0,0,170,250),(0,140,170,250),(0,198,170,250),(0,71,170,250),(177,71,170,250),(177,55,170,250),(177,55,180,250),(177,16,180,250),(177,16,180,14),(4,16,180,14),(230,16,180,14),(193,0,0,0),(0,39,0,0),(0,90,0,0),(0,221,0,0),(0,221,0,236),(36,221,0,236),(36,221,147,236),(36,221,147,73),(254,221,147,73),(254,221,197,73),(254,221,197,15),(254,182,197,15),(103,182,197,15),(163,182,197,15),(163,126,197,15),(163,181,197,15),(163,181,197,30),(163,7,197,30),(163,7,197,119),(13,7,197,119),(13,7,197,46),(13,7,197,190),(13,7,64,190),(13,7,64,166),(27,7,64,166),(0,0,55,0),(0,0,55,220),(198,0,55,220),(0,0,0,125),(188,0,0,125),(192,0,0,125),(192,0,0,102),(192,0,0,15),(192,248,0,15),(93,248,0,15),(93,248,164,15),(93,248,155,15),(73,248,155,15),(156,248,155,15),(156,248,155,183),(156,248,155,232),(156,248,155,79),(27,248,155,79),(27,248,155,73),(39,248,155,73),(39,248,155,84),(39,248,185,84),(39,248,229,84),(39,138,229,84),(39,138,16,84),(0,84,0,0),(121,84,0,0),(121,84,253,0),(121,84,253,49),(121,84,253,127),(121,84,222,127),(204,84,222,127),(204,84,87,127),(204,84,87,68),(0,0,0,114),(0,0,146,114),(0,0,146,130),(0,192,146,130),(0,71,146,130),(137,71,146,130),(137,5,146,130),(137,95,146,130),(137,95,146,183),(7,95,146,183),(7,95,71,183),(7,93,71,183),(22,93,71,183),(157,93,71,183),(157,93,71,60),(1,0,0,0),(1,0,170,0),(204,0,0,0),(204,0,0,171),(204,0,14,171),(64,0,14,171),(64,0,125,171),(64,0,226,171),(64,51,226,171),(251,51,226,171),(48,0,0,0),(66,0,0,0),(66,56,0,0),(66,56,174,0),(0,0,0,223),(0,32,0,223),(0,32,0,49),(0,185,0,0),(42,185,0,0),(72,185,0,0),(72,185,167,0),(118,185,167,0),(118,185,167,231),(243,185,167,231),(243,185,167,42),(243,185,167,29),(243,185,110,29),(123,185,110,29),(123,33,110,29),(43,33,110,29),(57,33,110,29),(57,33,110,233),(213,33,110,233),(213,33,110,151),(98,0,0,0),(68,0,0,0),(71,0,0,0),(71,0,0,102),(71,0,0,181),(71,0,143,181),(181,0,143,181),(181,0,81,181),(181,0,112,181),(181,51,112,181),(190,51,112,181),(0,222,0,0),(0,120,0,0),(93,120,0,0),(93,20,0,0),(93,140,0,0),(93,252,0,0),(0,7,0,0),(0,7,42,0),(234,7,42,0),(234,7,71,0),(234,206,71,0),(133,206,71,0),(183,0,0,0),(183,100,0,0),(28,100,0,0),(28,100,202,0),(28,162,202,0),(28,122,202,0),(103,122,202,0),(103,122,8,0),(118,122,8,0),(118,122,163,0),(140,122,163,0),(167,122,163,0),(167,122,75,0),(167,54,75,0),(73,54,75,0),(73,54,166,0),(104,54,166,0),(104,88,166,0),(0,0,0,203),(83,0,0,203),(83,120,0,203),(0,0,0,177),(152,0,0,177),(152,0,64,177),(152,77,64,177),(152,48,64,177),(74,48,64,177),(74,48,170,177),(202,48,170,177),(202,48,32,177),(202,48,202,177),(117,48,202,177),(12,48,202,177),(12,48,202,254),(12,48,202,70),(12,43,202,70),(247,43,202,70),(247,43,196,70),(247,43,137,70),(247,43,245,70),(247,43,245,120),(0,0,0,103),(0,0,45,103),(0,0,206,103),(0,169,206,103),(0,169,206,214),(0,169,206,71),(0,169,95,71),(0,169,95,212),(0,169,121,212),(0,0,0,88),(0,0,0,140),(0,0,0,40),(0,106,0,40),(0,106,0,113),(0,106,0,59),(0,106,225,59),(0,106,2,59),(0,106,2,55),(0,0,0,116),(229,0,0,116),(229,0,229,116),(229,0,68,116),(231,0,68,116),(126,0,68,116),(126,0,68,139),(126,0,68,205),(126,191,68,205),(126,191,68,246),(126,39,68,246),(126,39,68,90),(126,109,68,90),(126,109,68,98),(126,6,68,98),(11,6,68,98),(11,6,68,176),(11,164,68,176),(11,252,68,176),(11,170,68,176),(214,170,68,176),(214,170,234,176),(214,170,90,176),(0,0,199,0),(0,0,199,11),(0,0,202,11),(0,0,202,11),(0,0,202,214),(0,0,202,161),(0,80,202,161),(0,80,202,30),(0,112,202,30),(0,30,202,30),(0,30,202,67),(84,0,0,0),(84,251,0,0),(84,214,0,0),(84,202,0,0),(19,202,0,0),(19,56,0,0),(19,56,0,181),(19,73,0,181),(19,73,0,236),(19,29,0,236),(28,29,0,236),(28,29,0,27),(28,29,0,95),(28,29,0,244),(28,29,0,83),(28,29,0,213),(28,29,136,213),(27,29,136,213),(27,29,129,213),(0,0,0,66),(0,220,0,66),(66,220,0,66),(66,220,177,66),(66,220,177,17),(66,220,126,17),(168,220,126,17),(168,220,121,17),(168,220,64,17),(0,0,0,152),(48,0,0,152),(0,249,0,0),(0,249,69,0),(0,249,237,0),(0,249,237,53),(0,170,237,53),(0,170,237,30),(0,170,119,30),(0,0,146,0),(0,0,127,0),(0,0,161,0),(180,0,161,0),(180,0,110,0),(180,0,110,145),(180,131,110,145),(43,131,110,145),(43,131,165,145),(43,131,114,145),(43,129,114,145),(43,129,193,145),(43,129,193,240),(43,130,193,240),(43,130,193,8),(43,130,253,8),(43,130,253,86),(43,142,253,86),(0,9,0,0),(0,9,0,189),(76,0,0,0),(76,0,157,0),(76,42,157,0),(76,42,23,0),(76,42,93,0),(76,67,93,0),(88,67,93,0),(88,67,93,154),(119,67,93,154),(119,67,51,154),(0,148,0,0),(0,148,119,0),(0,0,0,217),(0,0,0,8),(0,0,0,92),(0,0,246,92),(0,0,160,92),(0,0,160,66),(0,2,160,66),(0,2,95,66),(0,244,95,66),(0,244,249,66),(0,244,69,66),(0,244,26,66),(0,244,92,66),(0,244,76,66),(0,244,173,66),(0,244,173,5),(0,244,254,5),(0,244,254,186),(158,244,254,186),(158,40,254,186),(158,40,225,186),(106,40,225,186),(106,40,225,188),(150,40,225,188),(150,252,225,188),(40,252,225,188),(40,252,225,146),(40,252,225,189),(0,75,0,0),(0,92,0,0),(0,92,88,0),(0,92,88,61),(176,92,88,61),(176,92,88,58),(148,92,88,58),(148,92,88,227),(148,171,88,227),(148,34,88,227),(175,34,88,227),(175,137,88,227),(175,212,88,227),(175,212,88,116),(175,212,213,116),(0,196,0,0),(0,132,0,0),(0,161,0,0),(0,161,89,0),(0,16,89,0),(0,16,89,179),(0,16,176,179),(45,16,176,179),(45,16,234,179),(45,16,234,239),(72,16,234,239),(219,16,234,239),(219,112,234,239),(219,112,212,239),(219,53,212,239),(219,53,231,239),(219,228,231,239),(219,228,231,117),(219,228,208,117),(219,228,208,167),(219,228,41,167),(51,228,41,167),(51,228,41,110),(0,0,67,0),(0,0,102,0),(0,97,102,0),(0,0,0,15),(166,0,0,15),(166,19,0,15),(221,19,0,15),(221,19,0,135),(67,19,0,135),(67,177,0,135),(116,177,0,135),(116,177,134,135),(116,177,219,135),(116,177,219,43),(116,177,219,158),(126,177,219,158),(126,168,219,158),(126,74,219,158),(0,165,0,0),(242,165,0,0),(176,165,0,0),(176,165,0,162),(224,165,0,162),(224,165,0,49),(224,165,34,49),(224,165,34,33),(224,165,126,33),(224,165,42,33),(0,0,0,20),(0,0,0,184),(64,0,0,184),(64,0,192,184),(64,0,51,184),(64,0,65,184),(64,0,65,155),(0,132,0,0),(0,132,216,0),(23,132,216,0),(23,132,216,56),(23,132,216,41),(23,132,165,41),(23,221,165,41),(23,87,165,41),(23,87,165,184),(23,23,165,184),(23,23,78,184),(23,23,78,199),(23,23,118,199),(135,23,118,199),(135,23,193,199),(135,23,193,82),(135,23,74,82),(135,23,21,82),(71,23,21,82),(71,23,21,139),(169,23,21,139),(169,23,21,76),(0,0,1,0),(0,152,1,0),(0,152,242,0),(0,152,27,0),(0,152,189,0),(0,152,8,0),(0,152,8,191),(0,152,8,242),(0,152,215,242),(0,152,122,242),(0,152,221,242),(0,233,221,242),(0,233,107,242),(0,233,190,242),(0,233,190,228),(142,233,190,228),(0,0,67,0),(0,214,67,0),(0,2,67,0),(34,2,67,0),(30,0,0,0),(30,0,216,0),(30,0,216,94),(120,0,216,94),(120,143,216,94),(221,143,216,94),(69,143,216,94),(215,143,216,94),(230,143,216,94),(0,0,0,12),(166,0,0,12),(141,0,0,12),(108,0,0,12),(108,0,0,234),(108,0,27,234),(108,0,190,234),(108,255,190,234),(108,255,101,234),(108,255,147,234),(108,10,147,234),(108,10,39,234),(108,10,39,219),(108,10,39,101),(0,0,253,0),(0,0,94,0),(0,0,244,0),(0,0,244,150),(0,0,244,132),(0,131,244,132),(0,131,244,21),(0,0,0,123),(0,7,0,123),(166,0,0,0),(166,72,0,0),(166,72,0,160),(59,72,0,160),(59,247,0,160),(59,247,120,160),(59,247,18,160),(59,247,132,160),(59,247,132,84),(59,36,132,84),(169,36,132,84),(169,36,8,84),(169,36,8,80),(169,36,8,222),(169,213,8,222),(169,213,8,246),(28,213,8,246),(63,213,8,246),(239,213,8,246),(239,213,8,176),(189,213,8,176),(24,213,8,176),(219,213,8,176),(219,213,8,201),(219,213,210,201),(18,213,210,201),(18,209,210,201),(18,209,210,95),(18,209,161,95),(111,209,161,95),(111,209,161,198),(111,200,161,198),(111,200,80,198),(111,200,198,198),(111,200,104,198),(0,0,121,0),(221,0,121,0),(221,0,121,130),(221,0,49,130),(221,0,49,11),(221,178,49,11),(221,178,19,11),(91,178,19,11),(0,0,0,252),(0,0,0,224),(0,0,68,224),(87,0,68,224),(87,0,112,224),(87,0,112,175),(87,0,112,22),(173,0,112,22),(173,0,215,22),(17,0,215,22),(17,0,215,10),(17,82,215,10),(17,82,216,10),(17,181,216,10),(130,181,216,10),(130,181,131,10),(130,181,131,144),(130,113,131,144),(229,0,0,0),(111,0,0,0),(111,0,40,0),(111,0,84,0),(165,0,84,0),(165,0,141,0),(78,0,141,0),(144,0,141,0),(0,0,0,50),(0,0,0,250),(0,0,0,164),(0,0,0,38),(0,0,0,137),(0,0,170,137),(0,0,170,206),(221,0,170,206),(221,111,170,206),(221,135,170,206),(252,135,170,206),(252,135,170,10),(58,135,170,10),(26,135,170,10),(63,135,170,10),(63,24,170,10),(63,35,170,10),(82,35,170,10),(123,35,170,10),(123,35,170,201),(123,35,170,240),(123,35,170,125),(123,35,170,103),(0,0,0,236),(0,122,0,236),(52,122,0,236),(52,239,0,236),(52,239,0,102),(92,239,0,102),(248,239,0,102),(185,239,0,102),(175,239,0,102),(0,0,0,159),(0,0,0,185),(27,0,0,185),(27,0,0,249),(27,0,21,249),(27,0,21,125),(27,0,95,125),(10,0,95,125),(10,81,95,125),(172,81,95,125),(172,165,95,125),(172,232,95,125),(96,0,0,0),(83,0,0,0),(83,73,0,0),(83,73,191,0),(83,73,121,0),(83,73,30,0),(83,73,30,227),(83,73,30,137),(152,73,30,137),(152,187,30,137),(152,187,30,112),(0,0,67,0),(0,0,212,0),(153,0,212,0),(81,0,212,0),(81,0,212,231),(236,0,0,0),(236,0,0,100),(236,0,0,154),(0,59,0,0),(0,59,15,0),(0,235,15,0),(23,235,15,0),(82,235,15,0),(30,235,15,0),(30,12,15,0),(0,158,0,0),(0,158,49,0),(0,158,49,165),(125,158,49,165),(125,158,49,187),(125,158,49,35),(125,158,95,35),(201,158,95,35),(189,158,95,35),(189,158,95,55),(0,0,0,130),(0,0,0,248),(0,0,137,248),(0,95,137,248),(0,121,137,248),(115,121,137,248),(0,0,62,0),(0,0,62,129),(0,0,62,218),(64,0,62,218),(167,0,62,218),(167,0,85,218),(167,0,85,110),(167,0,235,110),(167,0,235,80),(167,0,180,80),(167,0,180,149),(167,0,180,170),(167,233,180,170),(167,233,138,170),(167,244,138,170),(180,244,138,170),(180,27,138,170),(146,0,0,0),(146,0,0,165),(146,0,0,85),(26,0,0,85),(26,0,106,85),(26,89,106,85),(26,89,106,220),(26,89,106,171),(26,89,251,171),(26,158,251,171),(148,158,251,171),(24,158,251,171),(24,158,20,171),(65,158,20,171),(65,158,154,171),(65,158,63,171),(95,158,63,171),(95,158,70,171),(95,42,70,171),(95,42,70,206),(95,42,77,206),(95,42,77,217),(95,141,77,217),(95,119,77,217),(95,227,77,217),(95,39,77,217),(95,28,77,217),(95,28,142,217),(95,28,37,217),(127,28,37,217),(127,28,37,251),(0,0,191,0),(0,0,191,68),(0,122,191,68),(159,122,191,68),(159,122,238,68),(1,122,238,68),(61,122,238,68),(61,122,6,68),(61,122,6,31),(61,122,6,187),(125,122,6,187),(183,0,0,0),(183,0,0,155),(82,0,0,155),(82,29,0,155),(0,0,0,239),(0,0,0,243),(244,0,0,243),(244,171,0,243),(244,171,0,191),(244,171,223,191),(244,173,223,191),(244,173,223,208),(225,173,223,208),(225,173,223,183),(225,92,223,183),(35,92,223,183),(35,141,223,183),(35,193,223,183),(35,49,223,183),(35,231,223,183),(35,97,223,183),(0,0,117,0),(0,190,117,0),(0,190,22,0),(221,190,22,0),(221,190,142,0),(221,190,231,0),(0,14,0,0),(0,14,157,0),(124,14,157,0),(124,14,157,175),(124,14,157,44),(124,14,121,44),(124,14,121,204),(124,14,232,204),(67,14,232,204),(67,14,232,111),(67,14,21,111),(193,14,21,111),(0,0,39,0),(0,0,195,0),(0,194,195,0),(0,194,195,84),(0,194,195,44),(0,194,130,44),(0,194,135,44),(0,162,135,44),(0,181,135,44),(0,242,0,0),(0,0,239,0),(0,158,239,0),(0,131,239,0),(131,131,239,0),(0,72,0,0),(0,72,45,0),(229,0,0,0),(33,0,0,0),(33,0,22,0),(187,0,22,0),(37,0,22,0),(37,40,22,0),(37,40,22,237),(37,8,22,237),(37,8,22,217),(37,18,22,217),(37,80,22,217),(37,80,22,124),(214,80,22,124),(214,80,44,124),(58,0,0,0),(58,0,0,72),(58,0,147,72),(58,0,147,72),(214,0,147,72),(35,0,147,72),(37,0,147,72),(0,100,0,0),(0,100,0,240),(0,100,0,136),(0,100,190,136),(0,121,190,136),(0,121,40,136),(0,121,3,136),(0,121,3,88),(0,121,229,88),(0,121,229,172),(0,10,0,0),(0,142,0,0),(0,182,0,0),(0,73,0,0),(0,73,37,0),(0,19,0,0),(114,19,0,0),(114,19,0,34),(12,19,0,34),(12,226,0,34),(12,118,0,34),(12,118,0,104),(138,118,0,104),(138,118,0,116),(138,118,0,3),(138,190,0,3),(138,190,187,3),(138,190,187,198),(125,190,187,198),(0,217,0,0),(0,217,205,0),(0,126,205,0),(0,126,205,171),(0,4,205,171),(84,4,205,171),(211,4,205,171),(180,4,205,171),(78,4,205,171),(78,4,48,171),(0,206,0,0),(0,206,0,123),(0,206,0,87),(0,206,0,104),(0,0,180,0),(0,0,206,0),(0,0,240,0),(197,0,240,0),(197,173,240,0),(197,62,240,0),(197,241,240,0),(197,241,78,0),(197,241,78,78),(197,241,78,76),(197,35,78,76),(235,0,0,0),(195,0,0,0),(195,0,0,216),(195,0,0,3),(195,0,113,3),(195,184,113,3),(195,184,113,149),(195,147,113,149),(195,149,113,149),(0,201,0,0),(0,201,78,0),(0,254,78,0),(0,254,78,60),(214,254,78,60),(214,254,78,7),(214,254,78,211),(156,254,78,211),(156,254,153,211),(156,254,153,7),(156,123,153,7),(83,123,153,7),(83,123,153,247),(83,123,153,251),(83,123,153,232),(83,123,210,232),(152,123,210,232),(152,123,210,233),(27,123,210,233),(27,123,253,233),(27,123,253,215),(27,171,253,215),(27,171,13,215),(192,0,0,0),(192,0,0,222),(98,0,0,222),(45,0,0,222),(45,0,0,200),(0,0,0,159),(0,0,233,159),(0,196,0,0),(0,196,0,92),(179,196,0,92),(179,196,50,92),(153,196,50,92),(153,196,50,166),(153,196,50,140),(153,177,50,140),(153,177,154,140),(153,177,154,121),(153,177,186,121),(153,177,186,70),(153,62,186,70),(98,62,186,70),(240,0,0,0),(240,0,143,0),(68,0,143,0),(68,71,143,0),(229,71,143,0),(213,71,143,0),(213,248,143,0),(140,248,143,0),(140,49,143,0),(140,49,143,237),(140,49,25,237),(0,0,35,0),(0,207,35,0),(0,118,0,0),(0,118,0,144),(0,118,0,173),(0,118,0,104),(0,118,200,104),(0,118,200,88),(0,118,200,208),(200,118,200,208),(200,118,24,208),(200,118,4,208),(107,118,4,208),(107,172,4,208),(107,64,4,208),(107,64,196,208),(107,64,196,62),(77,64,196,62),(77,64,17,62),(77,64,132,62),(77,43,132,62),(77,127,132,62),(43,127,132,62),(43,127,132,147),(43,127,115,147),(58,127,115,147),(58,203,115,147),(138,203,115,147),(138,242,115,147),(138,242,130,147),(149,0,0,0),(175,0,0,0),(175,34,0,0),(175,238,0,0),(175,226,0,0),(175,224,0,0),(166,224,0,0),(166,151,0,0),(166,67,0,0),(166,67,35,0),(166,67,55,0),(166,67,100,0),(207,67,100,0),(190,67,100,0),(190,67,244,0),(190,67,255,0),(190,140,255,0),(190,183,255,0),(190,177,255,0),(133,177,255,0),(133,177,255,247),(9,177,255,247),(9,93,255,247),(9,51,255,247),(81,51,255,247),(81,216,255,247),(81,216,53,247),(105,216,53,247),(153,216,53,247),(153,216,53,79),(0,0,45,0),(0,0,45,123),(0,0,94,123),(0,0,34,123),(0,0,233,123),(120,0,233,123),(0,33,0,0),(0,33,211,0),(227,33,211,0),(227,66,211,0),(227,66,219,0),(0,0,79,0),(115,0,79,0),(115,0,79,35),(115,0,79,131),(73,0,79,131),(73,0,101,131),(200,0,101,131),(200,0,101,202),(200,221,101,202),(200,221,183,202),(141,221,183,202),(0,0,45,0),(0,0,45,51),(0,166,45,51),(100,166,45,51),(100,166,45,233),(141,166,45,233),(141,82,45,233),(141,82,45,26),(141,82,221,26),(55,82,221,26),(55,82,221,142),(55,82,125,142),(55,82,199,142),(41,82,199,142),(41,14,199,142),(114,14,199,142),(114,14,39,142),(114,6,39,142),(114,6,244,142),(114,6,201,142),(47,6,201,142),(47,6,230,142),(47,6,230,41),(47,6,230,150),(254,6,230,150),(254,6,157,150),(254,6,157,63),(254,6,157,225),(254,194,157,225),(254,194,25,225),(198,194,25,225),(198,29,25,225),(33,29,25,225),(33,29,65,225),(194,29,65,225),(194,29,65,54),(137,29,65,54),(137,67,65,54),(137,227,65,54),(35,0,0,0),(35,1,0,0),(209,1,0,0),(191,1,0,0),(184,1,0,0),(184,1,0,119),(103,1,0,119),(89,1,0,119),(89,1,0,38),(244,1,0,38),(148,0,0,0),(148,0,0,174),(32,0,0,174),(32,0,0,199),(0,0,228,0),(0,0,228,194),(0,14,228,194),(0,128,228,194),(232,128,228,194),(232,128,253,194),(232,128,253,212),(232,128,191,212),(232,128,201,212),(232,128,197,212),(0,0,0,92),(239,0,0,92),(239,131,0,92),(239,14,0,92),(84,14,0,92),(7,14,0,92),(0,193,0,0),(0,116,0,0),(0,116,51,0),(0,116,45,0),(0,116,45,136),(34,116,45,136),(0,46,0,0),(0,46,0,151),(0,46,223,151),(208,46,223,151),(208,46,223,80),(208,228,223,80),(208,228,223,9),(208,228,105,9),(208,252,105,9),(208,252,230,9),(208,252,126,9),(208,252,106,9),(208,52,106,9),(208,52,53,9),(208,52,53,112),(208,221,53,112),(208,221,53,156),(208,221,98,156),(154,221,98,156),(154,60,98,156),(154,60,34,156),(154,142,34,156),(154,208,34,156),(154,103,34,156),(110,103,34,156),(219,103,34,156),(219,103,129,156),(15,103,129,156),(51,103,129,156),(51,103,129,214),(51,103,129,219),(241,103,129,219),(241,103,169,219),(0,0,0,210),(0,0,168,210),(0,0,255,0),(0,0,0,65),(126,0,0,65),(186,0,0,65),(186,103,0,65),(186,31,0,65),(163,31,0,65),(163,31,182,65),(163,186,182,65),(205,186,182,65),(205,186,182,246),(172,186,182,246),(85,186,182,246),(85,186,206,246),(85,186,206,222),(85,186,255,222),(11,186,255,222),(11,186,255,173),(11,186,151,173),(11,186,151,151),(11,186,169,151),(11,186,169,183),(97,186,169,183),(97,186,63,183),(110,0,0,0),(110,250,0,0),(109,250,0,0),(65,0,0,0),(30,0,0,0),(147,0,0,0),(147,0,199,0),(147,0,199,199),(156,0,199,199),(156,0,99,199),(156,173,99,199),(156,173,99,205),(156,173,99,141),(156,30,99,141),(113,30,99,141),(113,30,177,141),(32,30,177,141),(192,30,177,141),(192,30,187,141),(192,119,187,141),(192,18,187,141),(192,205,187,141),(76,205,187,141),(76,159,187,141),(76,159,221,141),(219,159,221,141),(1,159,221,141),(1,84,221,141),(1,101,221,141),(234,101,221,141),(156,101,221,141),(156,101,128,141),(156,174,128,141),(156,212,128,141),(156,212,128,232),(156,44,128,232),(156,44,147,232),(156,44,147,53),(226,44,147,53),(78,44,147,53),(78,44,147,192),(78,44,147,77),(78,226,147,77),(78,226,146,77),(78,226,146,77),(78,226,87,77),(78,149,87,77),(78,149,24,77),(105,149,24,77),(105,149,151,77),(105,149,2,77),(0,0,83,0),(241,0,83,0),(241,220,83,0),(241,220,83,184),(241,220,98,184),(186,220,98,184),(186,220,148,184),(186,220,22,184),(186,220,22,169),(186,220,22,21),(139,0,0,0),(205,0,0,0),(205,135,0,0),(205,62,0,0),(205,62,152,0),(0,0,247,0),(0,0,247,99),(0,143,247,99),(100,143,247,99),(0,0,111,0),(224,0,111,0),(0,0,0,15),(0,74,0,15),(0,172,0,15),(0,172,146,15),(236,172,146,15),(236,154,146,15),(236,9,146,15),(236,9,146,109),(236,190,146,109),(236,88,146,109),(236,88,146,234),(236,88,52,234),(191,88,52,234),(139,88,52,234),(139,163,52,234),(139,163,124,234),(226,0,0,0),(226,0,232,0),(226,137,232,0),(226,137,232,56),(226,137,232,204),(226,119,232,204),(0,0,127,0),(0,0,131,0),(23,0,131,0),(23,0,125,0),(69,0,125,0),(69,48,125,0),(69,48,97,0),(69,48,153,0),(69,48,198,0),(69,48,198,220),(69,48,198,238),(190,48,198,238),(0,0,35,0),(15,0,35,0),(15,0,43,0),(15,184,43,0),(0,0,0,234),(0,51,0,234),(0,51,0,126),(0,51,28,126),(10,51,28,126),(169,51,28,126),(169,51,28,176),(169,51,84,176),(67,51,84,176),(67,51,174,176),(67,198,174,176),(67,198,174,127),(67,198,10,127),(67,198,149,127),(0,0,74,0),(0,194,74,0),(0,0,0,30),(0,0,0,241),(0,0,0,171),(0,0,0,233),(213,0,0,233),(213,0,119,233),(213,0,119,66),(213,0,53,66),(106,0,53,66),(67,0,53,66),(67,0,0,66),(67,119,0,66),(0,0,135,0),(0,128,135,0),(0,128,135,169),(222,128,135,169),(222,116,135,169),(136,116,135,169),(136,116,135,33),(170,116,135,33),(170,229,135,33),(82,229,135,33),(82,229,67,33),(255,229,67,33),(77,229,67,33),(77,229,133,33),(77,99,133,33),(77,238,133,33),(0,184,0,0),(0,184,0,74),(0,184,0,248),(0,184,0,137),(51,184,0,137),(51,184,0,24),(51,55,0,24),(51,66,0,24),(51,68,0,24),(51,109,0,24),(51,109,0,184),(51,109,73,184),(0,0,0,185),(0,127,0,185),(24,0,0,0),(49,0,0,0),(49,0,138,0),(49,0,138,52),(49,104,138,52),(49,104,207,52),(49,34,207,52),(49,34,241,52),(189,34,241,52),(68,34,241,52),(68,34,228,52),(199,34,228,52),(199,34,181,52),(199,5,181,52),(199,5,181,71),(159,5,181,71),(159,5,181,176),(159,5,181,176),(150,5,181,176),(150,248,181,176),(150,248,181,68),(150,156,181,68),(102,0,0,0),(103,0,0,0),(103,39,0,0),(103,39,0,142),(0,0,0,1),(0,0,0,68),(197,0,0,68),(232,0,0,68),(232,0,155,68),(232,190,155,68),(232,28,155,68),(0,78,0,0),(0,105,0,0),(0,105,3,0),(0,144,3,0),(0,144,14,0),(0,144,16,0),(0,94,16,0),(0,0,0,5),(94,0,0,0),(244,0,0,0),(244,0,120,0),(44,0,120,0),(44,0,196,0),(162,0,196,0),(162,0,34,0),(162,0,44,0),(162,0,45,0),(162,76,45,0),(162,23,45,0),(162,23,14,0),(162,23,157,0),(162,209,157,0),(0,6,0,0),(0,6,0,113),(164,6,0,113),(72,6,0,113),(72,6,227,113),(72,6,46,113),(72,6,52,113),(72,6,92,113),(72,22,92,113),(89,22,92,113),(89,22,18,113),(89,183,18,113),(194,183,18,113),(44,0,0,0),(225,0,0,0),(125,0,0,0),(125,200,0,0),(125,24,0,0),(125,24,169,0),(125,251,169,0),(162,251,169,0),(162,253,169,0),(162,253,116,0),(162,204,116,0),(69,204,116,0),(69,204,116,58),(69,242,116,58),(69,242,105,58),(95,242,105,58),(131,0,0,0),(131,0,115,0),(245,0,115,0),(245,232,115,0),(245,232,115,210),(15,232,115,210),(200,232,115,210),(200,232,210,210),(200,13,210,210),(200,13,210,115),(200,54,210,115),(0,0,0,137),(0,0,176,137),(0,0,170,137),(0,0,153,137),(0,0,153,80),(0,10,153,80),(0,10,162,80),(0,10,162,48),(35,10,162,48),(35,215,162,48),(35,215,152,48),(42,0,0,0),(42,0,0,218),(0,0,210,0),(0,0,210,79),(0,3,210,79),(39,3,210,79),(39,3,70,79),(39,197,70,79),(0,18,0,0),(99,18,0,0),(99,18,199,0),(99,100,199,0),(99,100,254,0),(99,95,254,0),(99,95,254,64),(182,95,254,64),(182,108,254,64),(182,108,254,147),(117,108,254,147),(117,100,254,147),(117,48,254,147),(117,48,119,147),(117,239,119,147),(117,239,224,147),(0,0,0,226),(219,0,0,226),(219,0,0,84),(219,250,0,84),(219,250,0,176),(21,250,0,176),(21,144,0,176),(58,144,0,176),(145,144,0,176),(145,144,0,45),(145,144,0,245),(145,144,0,232),(145,144,212,232),(145,87,212,232),(145,87,255,232),(145,87,255,223),(236,87,255,223),(236,59,255,223),(236,59,231,223),(181,59,231,223),(99,0,0,0),(99,205,0,0),(99,205,98,0),(85,205,98,0),(85,205,98,119),(85,205,21,119),(85,254,21,119),(85,254,21,207),(85,140,21,207),(85,140,21,200),(85,140,21,177),(85,140,21,24),(85,140,21,19),(85,27,21,19),(150,27,21,19),(150,27,227,19),(150,27,113,19),(150,27,204,19),(5,27,204,19),(5,27,204,23),(5,203,204,23),(5,203,133,23),(5,203,150,23),(5,120,150,23),(184,120,150,23),(184,120,150,140),(182,120,150,140),(0,0,57,0),(0,0,57,13),(0,0,60,13),(0,0,99,13),(137,0,99,13),(137,0,108,13),(43,0,108,13),(43,0,108,198),(216,0,108,198),(216,0,190,198),(216,0,151,198),(216,0,151,73),(216,0,239,73),(216,0,239,253),(216,0,172,253),(3,0,172,253),(3,0,144,253),(3,0,144,41),(72,0,144,41),(72,0,144,233),(105,0,144,233),(52,0,144,233),(52,149,144,233),(52,22,144,233),(196,22,144,233),(196,211,144,233),(0,0,0,156),(0,0,88,156),(64,0,88,156),(64,93,88,156),(64,229,88,156),(64,229,88,211),(179,229,88,211),(179,239,88,211),(223,239,88,211),(66,239,88,211),(66,239,88,90),(66,239,88,40),(66,239,64,40),(66,239,64,1),(66,172,64,1),(142,172,64,1),(142,172,96,1),(142,53,96,1),(142,53,60,1),(142,53,60,200),(142,31,60,200),(142,31,210,200),(142,31,210,29),(142,183,210,29),(142,189,210,29),(142,189,210,1),(142,46,210,1),(247,46,210,1),(247,46,248,1),(247,206,248,1),(247,70,248,1),(247,70,248,90),(247,70,248,88),(247,70,3,88),(247,70,208,88),(247,190,208,88),(247,190,208,183),(247,190,208,179),(247,190,208,94),(232,190,208,94),(232,190,208,144),(232,190,208,96),(232,160,208,96),(232,160,208,139),(232,150,208,139),(103,150,208,139),(196,150,208,139),(196,150,109,139),(0,0,0,139),(64,0,0,139),(0,0,43,0),(0,242,43,0),(2,242,43,0),(2,242,43,109),(221,242,43,109),(165,242,43,109),(165,242,43,110),(136,0,0,0),(136,0,78,0),(136,131,78,0),(136,117,78,0),(0,0,201,0),(0,0,87,0),(0,0,87,115),(0,236,87,115),(245,236,87,115),(245,236,13,115),(245,236,13,243),(73,236,13,243),(73,151,13,243),(73,156,13,243),(161,156,13,243),(161,195,13,243),(161,195,13,111),(249,195,13,111),(214,195,13,111),(214,195,13,212),(214,158,13,212),(214,158,0,212),(214,19,0,212),(214,19,0,225),(214,19,0,208),(214,19,0,79),(197,0,0,0),(0,0,0,202),(168,0,0,202),(61,0,0,202),(61,0,64,202),(61,0,64,234),(61,0,64,81),(61,132,64,81),(96,0,0,0),(96,0,0,76),(96,124,0,76),(0,0,0,140),(124,0,0,140),(124,0,122,140),(124,0,73,140),(53,0,73,140),(53,0,73,253),(53,0,66,253),(53,210,66,253),(53,210,66,46),(53,6,66,46),(53,6,234,46),(53,6,234,164),(53,6,234,85),(77,0,0,0),(77,142,0,0),(77,26,0,0),(77,26,0,142),(77,171,0,142),(77,171,96,142),(77,89,96,142),(77,89,178,142),(88,89,178,142),(68,89,178,142),(68,89,178,249),(68,89,178,78),(68,102,178,78),(68,102,95,78),(68,23,95,78),(68,26,95,78),(74,26,95,78),(74,26,95,127),(74,26,95,5),(74,26,95,144),(208,26,95,144),(208,118,95,144),(208,118,95,243),(208,118,236,243),(208,118,236,241),(181,118,236,241),(0,0,0,132),(0,238,0,132),(0,2,0,0),(180,2,0,0),(96,2,0,0),(96,85,0,0),(25,85,0,0),(30,0,0,0),(30,0,171,0),(30,0,171,159),(30,236,171,159),(16,236,171,159),(16,229,171,159),(138,229,171,159),(138,207,171,159),(138,154,171,159),(138,154,122,159),(138,154,152,159),(123,154,152,159),(253,154,152,159),(253,154,74,159),(253,154,199,159),(253,98,199,159),(253,142,199,159),(253,142,199,135),(253,142,73,135),(40,142,73,135),(190,142,73,135),(190,171,73,135),(190,220,73,135),(190,220,73,151),(190,220,73,73),(7,220,73,73),(7,172,73,73),(7,172,130,73),(7,35,130,73),(7,158,130,73),(7,158,219,73),(0,93,0,0),(0,93,0,143),(0,93,0,209),(0,93,128,209),(0,93,128,83),(0,93,128,76),(0,93,128,20),(0,93,83,20),(145,93,83,20),(145,93,12,20),(145,235,12,20),(145,235,82,20),(180,235,82,20),(123,235,82,20),(123,235,120,20),(123,126,120,20),(123,126,120,87),(123,126,237,87),(123,126,243,87),(123,126,243,205),(123,126,84,205),(123,126,84,144),(123,128,84,144),(97,128,84,144),(97,128,84,188),(97,128,229,188),(98,128,229,188),(98,171,229,188),(98,136,229,188),(98,85,229,188),(253,0,0,0),(116,0,0,0),(116,0,0,198),(116,230,0,198),(116,230,0,56),(116,230,0,118),(202,230,0,118),(91,230,0,118),(182,230,0,118),(30,230,0,118),(30,230,0,251),(30,230,214,251),(30,230,214,164),(30,230,128,164),(30,230,128,105),(30,230,128,181),(212,230,128,181),(184,230,128,181),(184,253,128,181),(184,253,173,181),(184,253,173,121),(0,0,106,0),(0,0,106,190),(0,68,106,190),(0,68,94,190),(0,100,94,190),(0,0,94,190),(0,0,94,142),(0,0,94,167),(117,0,94,167),(117,0,94,5),(117,0,245,5),(117,0,245,34),(61,0,245,34),(61,140,245,34),(46,140,245,34),(46,140,182,34),(46,247,182,34),(46,33,182,34),(46,43,182,34),(0,0,0,115),(0,0,251,115),(0,117,251,115),(0,117,160,115),(145,117,160,115),(145,117,108,115),(145,159,108,115),(0,0,0,196),(0,73,0,196),(0,73,147,196),(0,243,147,196),(0,0,0,0),(62,0,0,0),(62,0,92,0),(185,0,0,0),(185,0,0,177),(203,0,0,177),(5,0,0,177),(5,0,0,122),(169,0,0,122),(169,0,0,125),(169,0,201,125),(169,0,201,29),(169,0,201,66),(0,243,0,0),(0,225,0,0),(233,225,0,0),(233,225,0,48),(87,225,0,48),(87,225,0,45),(87,225,101,45),(165,225,101,45),(165,225,217,45),(173,225,217,45),(253,225,217,45),(253,225,15,45),(0,113,0,0),(0,237,0,0),(0,237,0,243),(0,237,0,76),(0,237,17,76),(0,96,17,76),(0,96,114,76),(0,213,114,76),(0,117,114,76),(0,117,174,76),(0,117,174,240),(0,107,174,240),(0,107,46,240),(0,107,46,247),(0,107,46,56),(0,107,46,121),(0,22,46,121),(0,208,46,121),(0,208,97,121),(7,208,97,121),(0,0,0,242),(0,0,190,242),(0,0,63,242),(0,210,63,242),(0,209,63,242),(0,165,63,242),(204,165,63,242),(204,59,63,242),(204,59,63,234),(204,59,63,232),(207,59,63,232),(207,59,219,232),(207,59,2,232),(207,59,168,232),(218,59,168,232),(218,59,168,249),(218,59,35,249),(12,59,35,249),(12,59,35,57),(12,58,35,57),(222,58,35,57),(222,58,122,57),(222,58,122,1),(222,58,170,1),(0,0,0,223),(157,0,0,223),(157,143,0,223),(157,143,0,188),(157,143,0,138),(157,143,192,138),(218,143,192,138),(218,143,174,138),(0,146,0,0),(0,146,0,219),(0,146,0,170),(0,240,0,170),(0,20,0,170),(0,20,88,170),(0,238,88,170),(0,238,25,170),(0,238,25,13),(117,238,25,13),(117,238,25,9),(117,230,25,9),(119,230,25,9),(214,230,25,9),(214,230,124,9),(0,208,0,0),(0,208,0,248),(20,208,0,248),(20,208,0,22),(20,208,0,55),(20,208,229,55),(20,208,229,58),(20,208,172,58),(20,208,16,58),(0,0,0,23),(0,0,10,23),(0,0,10,130),(173,0,10,130),(173,183,10,130),(173,183,10,84),(173,183,220,84),(212,0,0,0),(212,0,0,10),(212,0,0,189),(212,173,0,189),(212,18,0,189),(212,18,76,189),(0,0,0,155),(0,0,0,126),(0,150,0,126),(212,150,0,126),(212,230,0,126),(212,230,158,126),(36,230,158,126),(36,230,158,29),(36,164,158,29),(132,164,158,29),(49,164,158,29),(0,84,0,0),(114,84,0,0),(114,84,187,0),(0,0,0,251),(0,0,0,42),(146,0,0,0),(146,0,181,0),(207,0,181,0),(0,217,0,0),(121,217,0,0),(163,217,0,0),(163,217,0,244),(163,16,0,244),(163,16,0,166),(65,16,0,166),(65,16,224,166),(0,99,0,0),(0,99,0,76),(0,99,69,76),(0,99,69,177),(0,254,69,177),(204,254,69,177),(4,0,0,0),(4,0,0,166),(4,0,158,166),(4,0,158,39),(4,0,158,39),(4,0,49,39),(0,0,83,0),(0,0,83,17),(225,0,83,17),(225,96,83,17),(225,96,24,17),(34,0,0,0),(34,0,0,31),(34,109,0,31),(34,109,252,31),(79,109,252,31),(79,109,184,31),(79,109,184,35),(55,109,184,35),(55,109,184,19),(55,109,184,36),(55,109,218,36),(55,109,218,114),(55,109,218,218),(55,109,218,29),(55,109,25,29),(52,109,25,29),(52,109,25,73),(52,109,25,241),(52,109,65,241),(52,109,65,188),(86,109,65,188),(160,109,65,188),(41,109,65,188),(41,5,65,188),(41,5,232,188),(41,5,95,188),(10,5,95,188),(10,5,31,188),(113,5,31,188),(44,5,31,188),(44,5,18,188),(8,5,18,188),(0,0,0,160),(0,0,83,160),(12,0,83,160),(186,0,83,160),(0,0,161,0),(0,0,161,102),(0,0,143,102),(10,0,143,102),(10,241,143,102),(10,241,143,52),(10,241,184,52),(0,124,0,0),(0,124,64,0),(0,124,64,174),(0,124,64,129),(0,66,64,129),(38,66,64,129),(210,66,64,129),(117,66,64,129),(117,66,64,122),(0,40,0,0),(155,40,0,0),(8,0,0,0),(8,0,0,209),(162,0,0,209),(162,0,0,197),(0,122,0,0),(0,10,0,0),(168,10,0,0),(208,10,0,0),(208,10,221,0),(208,10,147,0),(208,10,147,82),(208,137,147,82),(63,137,147,82),(101,137,147,82),(101,155,147,82),(254,155,147,82),(254,155,147,222),(0,0,123,0),(0,45,123,0),(0,45,39,0),(0,45,39,98),(0,45,39,19),(0,45,165,19),(0,47,165,19),(0,125,165,19),(0,182,165,19),(0,24,0,0),(0,24,0,68),(0,24,82,68),(0,7,82,68),(255,7,82,68),(255,7,82,90),(255,7,82,208),(255,224,82,208),(29,224,82,208),(29,224,82,6),(29,216,82,6),(29,216,52,6),(29,38,52,6),(29,38,229,6),(137,38,229,6),(137,38,229,59),(137,38,229,45),(0,0,0,160),(0,40,0,160),(112,40,0,160),(112,40,0,191),(112,40,0,254),(112,40,0,1),(158,40,0,1),(158,18,0,1),(158,18,0,113),(0,0,25,0),(0,0,25,174),(0,184,25,174),(0,172,25,174),(0,172,25,44),(29,172,25,44),(162,172,25,44),(108,172,25,44),(108,172,25,128),(108,152,25,128),(108,214,25,128),(108,214,181,128),(108,214,24,128),(108,164,24,128),(108,164,18,128),(108,106,18,128),(36,106,18,128),(70,106,18,128),(70,106,246,128),(87,0,0,0),(87,0,0,190),(163,0,0,190),(0,135,0,0),(0,135,62,0),(0,135,150,0),(0,135,172,0),(0,135,6,0),(0,135,119,0),(199,135,119,0),(195,135,119,0),(195,135,119,67),(195,250,119,67),(195,250,119,79),(195,97,119,79),(195,97,119,163),(195,71,119,163),(195,177,119,163),(115,177,119,163),(115,84,119,163),(115,84,119,23),(115,84,119,231),(115,84,80,231),(115,160,80,231),(105,160,80,231),(60,0,0,0),(60,0,0,135),(60,0,120,135),(184,0,120,135),(184,0,81,135),(184,0,45,135),(67,0,45,135),(67,0,45,135),(68,0,45,135),(127,0,0,0),(127,128,0,0),(127,128,251,0),(127,128,0,0),(127,128,0,75),(127,128,174,75),(127,128,17,75),(127,167,17,75),(127,167,68,75),(127,239,68,75),(127,239,68,238),(127,99,68,238),(127,220,68,238),(127,220,10,238),(127,220,38,238),(127,220,38,193),(32,0,0,0),(168,0,0,0),(84,0,0,0),(84,0,0,213),(84,228,0,213),(84,132,0,213),(84,132,238,213),(194,132,238,213),(0,0,0,200),(0,0,58,200),(0,146,58,200),(0,146,58,203),(0,192,58,203),(0,0,162,0),(0,244,162,0),(0,244,162,248),(0,238,162,248),(0,238,117,248),(182,238,117,248),(122,238,117,248),(0,55,0,0),(105,55,0,0),(105,182,0,0),(105,182,0,234),(105,182,101,234),(105,182,144,234),(105,182,204,234),(105,182,204,138),(105,182,204,92),(0,123,0,0),(0,123,128,0),(139,0,0,0),(159,0,0,0),(159,112,0,0),(159,112,8,0),(159,117,8,0),(159,117,8,4),(159,252,8,4),(20,252,8,4),(0,0,145,0),(147,0,145,0),(66,0,145,0),(172,0,145,0),(220,0,145,0),(0,18,0,0),(254,0,0,0),(165,0,0,0),(165,0,30,0),(246,0,0,0),(15,0,0,0),(66,0,0,0),(66,0,89,0),(66,0,89,125),(239,0,89,125),(6,0,0,0),(6,31,0,0),(9,31,0,0),(226,31,0,0),(52,31,0,0),(52,31,216,0),(52,31,216,111),(52,175,216,111),(52,175,77,111),(91,175,77,111),(91,175,207,111),(91,175,219,111),(91,175,219,19),(185,175,219,19),(185,175,219,209),(190,175,219,209),(190,246,219,209),(190,246,219,152),(0,0,53,0),(0,80,0,0),(0,41,0,0),(193,41,0,0),(59,41,0,0),(0,14,0,0),(0,25,0,0),(0,25,0,128),(0,25,207,128),(0,25,111,128),(169,25,111,128),(167,25,111,128),(167,139,111,128),(167,25,111,128),(167,25,111,86),(104,25,111,86),(104,25,111,42),(104,164,111,42),(218,164,111,42),(232,164,111,42),(232,164,190,42),(232,164,212,42),(131,164,212,42),(131,164,254,42),(131,164,254,42),(131,162,254,42),(131,27,254,42),(229,27,254,42),(27,27,254,42),(27,212,254,42),(27,212,254,152),(27,212,254,88),(27,212,254,234),(233,212,254,234),(233,212,92,234),(233,212,181,234),(233,195,181,234),(233,116,181,234),(233,116,181,238),(233,1,181,238),(233,1,181,57),(233,1,181,129),(233,1,171,129),(27,1,171,129),(14,1,171,129),(0,0,105,0),(0,0,105,56),(0,0,220,56),(0,243,220,56),(0,243,220,99),(2,243,220,99),(2,161,220,99),(34,161,220,99),(182,161,220,99),(182,161,220,164),(50,161,220,164),(22,161,220,164),(22,161,220,94),(22,161,220,88),(22,160,220,88),(157,160,220,88),(157,160,220,208),(157,69,220,208),(237,69,220,208),(237,69,220,166),(237,69,37,166),(237,69,37,145),(237,73,37,145),(53,0,0,0),(53,0,0,130),(222,0,0,130),(10,0,0,130),(10,0,150,130),(231,0,150,130),(234,0,150,130),(0,75,0,0),(0,75,0,15),(0,96,0,0),(0,96,142,0),(0,96,179,0),(54,96,179,0),(54,96,148,0),(54,96,171,0),(172,96,171,0),(172,96,157,0),(172,96,157,164),(172,96,115,164),(172,96,115,204),(216,96,115,204),(81,0,0,0),(81,0,32,0),(81,0,115,0),(81,0,71,0),(81,0,71,253),(81,0,40,253),(53,0,40,253),(116,0,40,253),(0,0,191,0),(134,0,191,0),(134,0,191,29),(134,0,191,235),(134,84,191,235),(134,84,162,235),(134,84,153,235),(134,84,240,235),(134,84,240,111),(134,34,240,111),(134,34,29,111),(134,34,29,166),(134,34,29,85),(245,34,29,85),(65,34,29,85),(65,252,29,85),(98,252,29,85),(98,123,29,85),(235,123,29,85),(235,87,29,85),(235,87,29,218),(235,219,29,218),(235,219,29,130),(198,219,29,130),(198,219,29,166),(198,163,29,166),(198,163,188,166),(198,163,203,166),(194,163,203,166),(194,163,194,166),(228,163,194,166),(0,55,0,0),(0,55,55,0),(0,55,67,0),(0,55,67,73),(0,55,67,222),(0,55,67,242),(0,55,67,249),(0,55,67,89),(0,55,67,114),(0,55,67,137),(0,55,67,231),(48,55,67,231),(48,77,67,231),(71,77,67,231),(71,219,67,231),(71,219,67,2),(82,219,67,2),(242,219,67,2),(242,219,74,2),(242,88,74,2),(242,88,3,2),(242,88,3,114),(218,88,3,114),(0,106,0,0),(0,106,13,0),(0,0,0,127),(0,0,0,185),(112,0,0,185),(112,208,0,185),(222,208,0,185),(113,0,0,0),(0,0,226,0),(0,0,226,51),(126,0,226,51),(126,14,226,51),(126,14,226,247),(126,14,157,247),(126,14,108,247),(126,241,108,247),(126,241,108,68),(126,241,200,68),(126,32,200,68),(126,32,207,68),(126,32,70,68),(126,32,70,232),(126,32,70,108),(126,32,218,108),(126,32,68,108),(21,32,68,108),(21,32,169,108),(21,84,169,108),(21,84,169,4),(21,84,142,4),(21,84,66,4),(21,208,66,4),(21,208,188,4),(21,208,188,0),(21,208,188,101),(21,208,188,129),(21,208,65,129),(21,208,135,129),(52,208,135,129),(52,208,135,108),(70,208,135,108),(151,208,135,108),(151,208,135,179),(59,208,135,179),(240,208,135,179),(240,208,135,114),(240,212,135,114),(240,212,135,158),(240,212,91,158),(122,212,91,158),(34,212,91,158),(34,212,217,158),(34,212,217,24),(34,255,217,24),(34,255,217,126),(34,255,253,126),(34,167,253,126),(34,167,246,126),(107,167,246,126),(43,167,246,126),(43,167,246,71),(43,83,246,71),(43,83,145,71),(136,83,145,71),(136,83,2,71),(136,83,2,189),(120,83,2,189),(120,83,149,189),(120,41,149,189),(0,0,168,0),(0,0,168,29),(0,0,0,183),(0,167,0,183),(0,167,0,126),(0,90,0,126),(0,29,0,126),(0,0,0,13),(0,49,0,13),(0,0,0,16),(0,0,0,81),(0,0,153,81),(0,162,153,81),(116,162,153,81),(116,56,153,81),(116,56,153,153),(116,122,153,153),(128,122,153,153),(0,223,0,0),(0,0,0,133),(0,0,67,133),(150,0,67,133),(150,0,67,8),(150,0,72,8),(225,0,0,0),(225,0,122,0),(225,0,21,0),(225,0,21,154),(225,0,50,154),(225,0,16,154),(225,40,16,154),(225,40,159,154),(101,40,159,154),(79,40,159,154),(79,40,159,218),(96,40,159,218),(96,165,159,218),(96,165,145,218),(235,0,0,0),(235,0,0,157),(202,0,0,157),(202,242,0,157),(150,242,0,157),(150,242,0,175),(21,242,0,175),(21,242,47,175),(21,242,47,90),(21,242,83,90),(21,242,147,90),(21,242,147,243),(21,242,147,220),(21,242,147,11),(99,242,147,11),(166,242,147,11),(166,242,147,116),(134,242,147,116),(134,39,147,116),(134,39,76,116),(134,39,76,95),(134,39,165,95),(160,39,165,95),(160,39,165,201),(119,39,165,201),(119,39,165,0),(119,39,241,0),(127,0,0,0),(127,78,0,0),(224,78,0,0),(224,78,81,0),(224,124,81,0),(105,124,81,0),(105,124,81,66),(105,124,81,222),(0,0,144,0),(41,0,144,0),(0,0,21,0),(0,0,117,0),(0,0,117,15),(0,93,117,15),(0,158,117,15),(202,158,117,15),(202,158,72,15),(202,158,65,15),(202,238,65,15),(202,48,65,15),(202,160,65,15),(202,160,127,15),(202,181,127,15),(202,181,127,186),(0,163,0,0),(0,163,0,13),(62,163,0,13),(62,180,0,13),(0,0,0,47),(0,0,213,47),(0,0,213,36),(159,0,213,36),(0,0,43,0),(236,0,43,0),(90,0,43,0),(19,0,0,0),(19,0,22,0),(12,0,22,0),(12,0,22,252),(12,0,22,25),(12,15,22,25),(12,15,22,88),(0,251,0,0),(231,251,0,0),(133,251,0,0),(133,251,221,0),(133,251,84,0),(133,43,84,0),(133,58,84,0),(133,157,84,0),(133,157,30,0),(133,157,157,0),(133,157,49,0),(133,127,49,0),(141,127,49,0),(0,0,68,0),(0,39,68,0),(13,39,68,0),(252,39,68,0),(252,39,38,0),(252,157,38,0),(0,182,0,0),(0,182,172,0),(0,182,172,102),(0,182,213,102),(0,182,213,36),(0,182,213,78),(144,182,213,78),(0,52,0,0),(0,204,0,0),(188,0,0,0),(188,0,59,0),(188,0,59,113),(232,0,59,113),(232,83,59,113),(232,236,59,113),(178,236,59,113),(178,236,135,113),(178,193,135,113),(243,193,135,113),(243,193,135,132),(117,193,135,132),(117,193,156,132),(15,193,156,132),(63,193,156,132),(63,193,156,223),(63,193,52,223),(63,193,48,223),(205,193,48,223),(211,193,48,223),(244,193,48,223),(216,193,48,223),(205,193,48,223),(205,193,74,223),(205,193,20,223),(199,193,20,223),(199,15,20,223),(199,36,20,223),(199,36,70,223),(199,36,24,223),(199,121,24,223),(199,33,24,223),(199,125,24,223),(199,125,238,223),(238,125,238,223),(238,225,238,223),(238,225,121,223),(79,225,121,223),(79,225,121,33),(79,179,121,33),(79,179,121,210),(10,179,121,210),(10,179,51,210),(10,179,61,210),(10,179,61,113),(10,179,144,113),(44,0,0,0),(44,0,0,177),(44,0,114,177),(25,0,114,177),(25,196,114,177),(25,196,114,14),(25,196,116,14),(25,30,116,14),(77,30,116,14),(143,30,116,14),(143,174,116,14),(242,174,116,14),(242,174,116,47),(242,174,26,47),(242,174,26,81),(0,0,80,0),(0,0,80,116),(161,0,80,116),(161,0,80,98),(161,0,241,98),(161,0,241,36),(177,0,241,36),(177,0,92,36),(177,0,7,36),(177,0,51,36),(177,0,162,36),(177,0,101,36),(53,0,101,36),(53,9,101,36),(53,9,218,36),(53,9,218,178),(53,9,218,245),(53,9,218,213),(53,9,218,162),(53,9,218,56),(53,9,135,56),(164,9,135,56),(164,9,130,56),(164,45,130,56),(69,45,130,56),(72,45,130,56),(72,45,130,4),(31,45,130,4),(31,173,130,4),(25,173,130,4),(0,234,0,0),(0,234,0,202),(226,234,0,202),(226,156,0,202),(226,156,0,168),(226,75,0,168),(226,75,232,168),(172,75,232,168),(172,70,232,168),(152,70,232,168),(152,70,232,185),(0,0,165,0),(155,0,165,0),(0,0,166,0),(0,0,52,0),(0,0,52,88),(0,135,52,88),(216,135,52,88),(216,135,52,228),(216,135,149,228),(216,160,149,228),(216,160,152,228),(216,160,152,204),(216,160,152,30),(242,160,152,30),(242,37,152,30),(242,37,98,30),(242,184,98,30),(242,67,98,30),(242,67,12,30),(242,67,12,252),(60,67,12,252),(60,55,12,252),(60,55,63,252),(60,55,45,252),(60,55,155,252),(60,55,88,252),(60,55,88,12),(165,55,88,12),(165,100,88,12),(247,100,88,12),(247,100,88,204),(247,100,88,228),(247,100,88,52),(247,100,88,175),(247,218,88,175),(0,128,0,0),(0,128,0,230),(0,79,0,230),(0,80,0,230),(0,0,0,210),(0,172,0,210),(127,172,0,210),(40,172,0,210),(40,51,0,210),(0,168,0,0),(0,168,0,145),(0,168,60,145),(0,168,151,145),(0,168,252,145),(0,77,252,145),(49,0,0,0),(49,204,0,0),(49,204,206,0),(0,0,0,185),(0,0,0,228),(0,81,0,228),(0,81,0,243),(0,81,0,71),(5,81,0,71),(5,81,0,209),(5,81,220,209),(5,81,220,61),(5,81,82,61),(5,60,82,61),(5,171,82,61),(5,171,82,106),(5,171,82,1),(5,54,82,1),(5,222,82,1),(5,222,82,175),(240,222,82,175),(240,73,82,175),(164,73,82,175),(164,73,177,175),(164,73,172,175),(164,169,172,175),(155,169,172,175),(155,224,172,175),(155,115,172,175),(155,157,172,175),(0,208,0,0),(0,208,229,0),(0,14,229,0),(255,14,229,0),(171,14,229,0),(171,235,229,0),(173,235,229,0),(243,235,229,0),(50,235,229,0),(50,173,229,0),(50,173,229,195),(50,231,229,195),(50,231,31,195),(0,0,0,9),(0,0,0,108),(0,113,0,108),(0,97,0,108),(0,97,0,74),(191,97,0,74),(79,97,0,74),(79,49,0,74),(0,0,169,0),(0,0,78,0),(0,237,78,0),(0,237,64,0),(0,135,0,0),(0,135,94,0),(0,151,94,0),(129,151,94,0),(0,0,0,91),(0,193,0,91),(0,193,240,91),(0,193,240,49),(0,88,240,49),(0,138,240,49),(29,138,240,49),(0,0,0,174),(0,0,0,104),(0,0,219,0),(0,148,219,0),(0,46,219,0),(0,0,0,115),(60,0,0,115),(60,221,0,115),(0,232,0,0),(0,0,7,0),(0,0,7,235),(0,0,225,0),(0,40,225,0),(5,40,225,0),(5,40,144,0),(5,40,144,98),(5,40,144,36),(5,230,144,36),(5,230,144,156),(5,30,144,156),(252,0,0,0),(252,0,201,0),(12,0,201,0),(125,0,201,0),(125,0,171,0),(125,0,126,0),(125,5,126,0),(125,5,44,0),(127,5,44,0),(110,0,0,0),(110,208,0,0),(47,0,0,0),(47,0,0,222),(47,0,0,0),(47,0,0,37),(174,0,0,37),(174,0,0,80),(174,0,0,40),(0,0,222,0),(0,85,222,0),(0,195,222,0),(0,0,0,126),(0,0,76,126),(0,0,76,103),(0,0,76,175),(157,0,76,175),(151,0,76,175),(151,96,76,175),(151,96,167,175),(151,140,167,175),(164,0,0,0),(164,0,0,143),(164,0,0,219),(164,91,0,219),(164,53,0,219),(0,0,149,0),(0,0,24,0),(175,0,24,0),(175,220,24,0),(230,220,24,0),(230,220,238,0),(230,184,238,0),(127,184,238,0),(127,184,238,72),(0,0,46,0),(0,224,46,0),(0,249,46,0),(0,33,46,0),(0,33,127,0),(0,232,127,0),(0,232,127,183),(0,19,127,183),(0,16,127,183),(0,16,195,183),(0,16,195,172),(0,16,35,172),(142,16,35,172),(142,16,35,163),(0,0,221,0),(60,0,221,0),(60,0,221,252),(60,0,140,252),(60,0,140,120),(0,0,172,0),(0,0,226,0),(0,0,226,163),(119,0,226,163),(119,0,157,163),(119,0,18,163),(119,0,162,163),(98,0,162,163),(108,0,162,163),(108,0,68,163),(74,0,68,163),(177,0,68,163),(0,81,0,0),(245,81,0,0),(21,81,0,0),(21,81,0,142),(21,81,0,11),(17,81,0,11),(134,81,0,11),(134,81,29,11),(90,81,29,11),(154,81,29,11),(154,106,29,11),(154,106,170,11),(225,106,170,11),(225,231,170,11),(183,231,170,11),(206,0,0,0),(206,0,153,0),(254,0,153,0),(2,0,153,0),(2,0,192,0),(2,0,192,117),(173,0,192,117),(149,0,192,117),(149,2,192,117),(0,0,0,215),(0,0,0,30),(0,91,0,30),(60,91,0,30),(60,91,0,120),(200,91,0,120),(200,91,0,188),(200,207,0,188),(255,207,0,188),(255,207,0,55),(255,207,86,55),(255,207,86,106),(255,207,21,106),(150,207,21,106),(150,237,21,106),(150,237,21,209),(48,237,21,209),(45,237,21,209),(45,237,21,171),(189,237,21,171),(189,45,21,171),(189,253,21,171),(189,253,21,221),(189,47,21,221),(68,47,21,221),(68,162,21,221),(68,162,21,44),(68,162,251,44),(68,162,72,44),(68,162,72,178),(68,98,72,178),(186,98,72,178),(186,98,72,12),(61,98,72,12),(61,98,80,12),(61,98,247,12),(61,98,25,12),(61,160,25,12),(61,160,25,190),(61,175,25,190),(61,175,25,74),(61,175,25,49),(135,175,25,49),(135,175,49,49),(135,21,49,49),(37,21,49,49),(236,21,49,49),(236,21,164,49),(236,21,164,222),(236,21,107,222),(236,21,36,222),(236,212,36,222),(236,212,36,9),(104,212,36,9),(45,212,36,9),(45,212,43,9),(45,212,163,9),(45,147,163,9),(45,78,163,9),(45,78,76,9),(45,78,76,255),(45,181,76,255),(45,181,76,142),(45,217,76,142),(45,26,76,142),(45,26,30,142),(45,26,196,142),(45,26,196,151),(45,26,196,213),(35,26,196,213),(0,54,0,0),(0,0,94,0),(0,0,0,247),(195,0,0,247),(195,222,0,247),(195,222,0,43),(195,222,250,43),(195,222,164,43),(133,222,164,43),(133,210,164,43),(133,210,164,149),(61,210,164,149),(61,65,164,149),(61,65,164,106),(0,0,118,0),(32,0,118,0),(32,0,104,0),(32,109,104,0),(32,109,213,0),(32,109,213,170),(32,109,213,70),(32,109,167,70),(15,109,167,70),(15,109,236,70),(15,109,0,70),(15,109,76,70),(15,109,148,70),(15,149,148,70),(15,149,192,70),(15,149,63,70),(15,149,114,70),(0,93,0,0),(0,171,0,0),(0,171,168,0),(0,31,168,0),(0,31,210,0),(0,245,210,0),(0,68,210,0),(81,68,210,0),(96,68,210,0),(96,68,210,237),(209,68,210,237),(209,146,210,237),(71,146,210,237),(71,130,210,237),(0,0,213,0),(0,0,22,0),(0,189,22,0),(97,189,22,0),(97,189,22,37),(97,189,69,37),(97,239,69,37),(97,239,205,37),(236,239,205,37),(26,239,205,37),(26,127,205,37),(26,127,35,37),(26,127,227,37),(202,127,227,37),(202,53,227,37),(116,53,227,37),(3,53,227,37),(0,0,0,22),(0,0,0,204),(0,166,0,204),(170,166,0,204),(186,166,0,204),(186,166,112,204),(186,166,242,204),(193,166,242,204),(59,166,242,204),(59,166,242,53),(59,154,242,53),(59,33,242,53),(255,33,242,53),(53,33,242,53),(53,33,68,53),(53,33,68,92),(100,33,68,92),(0,0,142,0),(124,0,142,0),(124,250,142,0),(124,250,82,0),(124,181,82,0),(124,50,82,0),(124,16,82,0),(124,229,82,0),(124,229,139,0),(0,108,0,0),(0,173,0,0),(0,167,0,0),(0,167,0,198),(186,167,0,198),(11,167,0,198),(11,167,148,198),(11,167,93,198),(0,0,101,0),(0,51,101,0),(0,106,101,0),(202,106,101,0),(202,124,101,0),(202,124,99,0),(128,124,99,0),(0,0,0,134),(0,0,89,134),(73,0,89,134),(0,0,89,134),(0,128,89,134),(0,128,89,161),(126,128,89,161),(126,128,196,161),(126,128,22,161),(90,128,22,161),(90,128,22,181),(90,128,22,175),(0,175,0,0),(0,175,202,0),(0,175,41,0),(0,175,46,0),(0,175,46,90),(100,175,46,90),(100,175,46,71),(100,175,46,70),(100,175,108,70),(100,175,71,70),(248,175,71,70),(248,175,184,70),(2,175,184,70),(0,0,37,0),(0,118,37,0),(0,118,118,0),(0,118,88,0),(0,118,22,0),(64,118,22,0),(64,118,22,56),(64,118,164,56),(64,166,164,56),(64,146,164,56),(0,165,0,0),(0,165,0,219),(0,165,0,52),(0,145,0,52),(0,232,0,52),(0,111,0,52),(0,111,236,52),(0,111,9,52),(36,111,9,52),(36,220,9,52),(188,220,9,52),(188,220,9,144),(188,220,9,243),(188,220,142,243),(188,220,129,243),(188,220,129,151),(188,109,129,151),(188,11,129,151),(188,11,129,16),(188,11,129,213),(188,11,251,213),(188,14,251,213),(188,245,251,213),(188,245,150,213),(129,245,150,213),(129,245,102,213),(210,245,102,213),(210,245,238,213),(210,245,239,213),(210,245,239,29),(210,245,27,29),(210,245,27,211),(210,245,31,211),(210,223,31,211),(99,0,0,0),(99,0,57,0),(99,188,57,0),(225,188,57,0),(225,188,57,227),(225,188,57,115),(69,188,57,115),(69,188,57,30),(249,188,57,30),(249,110,57,30),(169,110,57,30),(0,0,0,175),(131,0,0,175),(131,0,0,48),(131,0,241,48),(0,87,0,0),(0,0,195,0),(0,125,195,0),(102,125,195,0),(102,80,195,0),(102,89,195,0),(102,89,26,0),(102,89,142,0),(102,35,142,0),(17,35,142,0),(17,35,37,0),(17,35,37,26),(17,8,37,26),(17,43,37,26),(17,43,37,195),(17,43,37,173),(17,43,37,30),(118,43,37,30),(118,43,51,30),(118,43,241,30),(118,199,241,30),(151,199,241,30),(0,0,0,34),(242,0,0,34),(0,0,221,0),(0,0,250,0),(0,253,250,0),(0,253,183,0),(0,205,183,0),(0,114,183,0),(0,186,183,0),(124,186,183,0),(124,186,86,0),(124,191,86,0),(174,191,86,0),(161,0,0,0),(161,0,0,190),(161,0,244,190),(161,0,244,114),(87,0,0,0),(45,0,0,0),(45,0,0,138),(45,0,150,138),(45,0,212,138),(45,0,156,138),(29,0,156,138),(0,0,0,193),(0,0,70,0),(0,217,70,0),(166,217,70,0),(166,217,70,254),(166,217,70,171),(113,217,70,171),(109,217,70,171),(109,217,125,171),(127,217,125,171),(191,217,125,171),(191,217,125,62),(191,29,125,62),(191,29,125,234),(191,29,108,234),(191,29,108,173),(191,29,108,131),(191,29,108,0),(191,7,108,0),(131,7,108,0),(131,7,22,0),(131,7,171,0),(232,7,171,0),(115,7,171,0),(115,247,171,0),(115,247,173,0),(115,247,173,246),(251,247,173,246),(251,247,183,246),(184,247,183,246),(184,247,183,169),(141,247,183,169),(141,191,183,169),(44,191,183,169),(232,191,183,169),(232,191,147,169),(215,191,147,169),(215,191,107,169),(215,125,107,169),(215,220,107,169),(0,0,0,235),(60,0,0,235),(0,59,0,0),(0,41,0,0),(230,41,0,0),(60,41,0,0),(173,41,0,0),(173,41,0,6),(173,154,0,6),(173,154,134,6),(208,154,134,6),(208,154,134,245),(208,154,134,72),(208,117,134,72),(208,117,134,217),(208,117,134,221),(205,0,0,0),(68,0,0,0),(68,0,206,0),(156,0,206,0),(245,0,206,0),(245,39,206,0),(109,39,206,0),(109,39,147,0),(109,39,43,0),(109,39,203,0),(109,20,203,0),(109,20,167,0),(109,20,189,0),(109,20,189,75),(109,223,189,75),(109,13,189,75),(175,13,189,75),(175,13,236,75),(175,252,236,75),(175,252,44,75),(55,252,44,75),(55,252,44,164),(55,252,56,164),(55,252,56,66),(55,252,173,66),(236,252,173,66),(125,252,173,66),(125,252,173,15),(125,252,173,103),(125,114,173,103),(0,0,229,0),(154,0,229,0),(154,0,71,0),(253,0,71,0),(0,220,0,0),(0,220,157,0),(180,220,157,0),(0,0,0,86),(0,0,214,86),(251,0,214,86),(251,210,214,86),(0,0,105,0),(0,0,105,244),(0,0,105,106),(0,0,105,167),(0,0,105,14),(0,186,105,14),(0,55,105,14),(0,55,55,14),(0,55,181,14),(0,166,181,14),(0,166,128,14),(0,121,128,14),(0,121,128,179),(0,121,110,179),(45,0,0,0),(45,0,0,31),(155,0,0,31),(155,248,0,31),(211,248,0,31),(211,248,55,31),(211,248,55,143),(211,248,55,112),(174,248,55,112),(253,248,55,112),(20,248,55,112),(120,248,55,112),(0,248,55,112),(0,248,135,112),(0,248,180,112),(0,248,96,112),(0,0,23,0),(0,0,5,0),(0,0,56,0),(0,58,56,0),(220,58,56,0),(220,58,56,209),(77,0,0,0),(77,146,0,0),(77,17,0,0),(77,17,173,0),(77,17,173,210),(77,17,224,210),(77,17,191,210),(77,17,205,210),(10,0,0,0),(196,0,0,0),(216,0,0,0),(0,0,172,0),(0,169,172,0),(214,169,172,0),(214,233,172,0),(214,233,181,0),(214,233,181,218),(214,208,181,218),(254,208,181,218),(254,200,181,218),(168,200,181,218),(168,200,181,139),(50,200,181,139),(50,200,24,139),(50,200,24,178),(50,200,24,193),(50,200,8,193),(50,200,7,193),(50,200,93,193),(196,200,93,193),(196,40,93,193),(152,0,0,0),(152,0,114,0),(152,0,114,186),(152,0,31,186),(152,0,31,41),(0,0,0,157),(177,0,0,157),(177,0,67,157),(177,90,67,157),(177,90,67,98),(177,90,54,98),(130,90,54,98),(130,241,54,98),(130,91,54,98),(130,91,54,121),(130,91,106,121),(130,91,106,61),(204,91,106,61),(204,91,100,61),(204,91,100,110),(204,232,100,110),(204,232,197,110),(204,51,197,110),(177,51,197,110),(177,21,197,110),(177,21,84,110),(177,21,155,110),(254,21,155,110),(254,130,155,110),(254,130,155,65),(254,130,100,65),(254,143,100,65),(254,143,29,65),(247,143,29,65),(247,128,29,65),(247,19,29,65),(247,19,82,65),(247,164,82,65),(177,164,82,65),(177,164,178,65),(177,164,178,209),(177,164,178,127),(190,164,178,127),(190,164,178,79),(190,164,5,79),(224,0,0,0),(52,0,0,0),(52,0,0,123),(52,0,88,123),(27,0,88,123),(27,0,88,29),(27,225,88,29),(71,225,88,29),(42,225,88,29),(42,225,88,184),(42,225,88,30),(42,206,88,30),(42,206,88,149),(42,182,88,149),(193,182,88,149),(193,182,214,149),(193,182,214,129),(0,138,0,0),(0,117,0,0),(10,117,0,0),(152,117,0,0),(152,117,55,0),(152,117,55,82),(152,117,55,245),(152,117,55,165),(239,117,55,165),(239,202,55,165),(239,202,209,165),(239,164,209,165),(239,215,209,165),(35,215,209,165),(35,55,209,165),(35,66,209,165),(35,66,120,165),(35,66,120,136),(0,0,89,0),(0,0,69,0),(0,0,69,237),(0,210,69,237),(0,179,69,237),(0,179,71,237),(0,0,71,237),(0,186,71,237),(87,186,71,237),(87,186,22,237),(87,186,22,56),(87,186,123,56),(254,186,123,56),(71,186,123,56),(71,57,123,56),(71,57,38,56),(0,0,150,0),(243,0,150,0),(243,0,177,0),(243,0,177,106),(243,0,104,106),(243,80,104,106),(217,80,104,106),(217,80,175,106),(204,80,175,106),(204,80,223,106),(204,80,223,102),(130,80,223,102),(130,72,223,102),(250,72,223,102),(146,72,223,102),(146,72,223,204),(206,0,0,0),(206,60,0,0),(0,184,0,0),(0,71,0,0),(0,118,0,0),(0,65,0,0),(0,65,156,0),(157,65,156,0),(72,65,156,0),(72,65,156,228),(72,200,156,228),(72,135,156,228),(27,0,0,0),(27,0,154,0),(24,0,154,0),(24,224,154,0),(160,224,154,0),(160,77,154,0),(160,77,100,0),(160,122,100,0),(160,122,201,0),(0,0,188,0),(0,178,188,0),(0,0,0,87),(0,0,5,87),(0,244,0,0),(0,248,0,0),(0,128,0,0),(0,172,0,0),(0,0,0,254),(74,0,0,254),(74,11,0,254),(74,190,0,254),(74,206,0,254),(73,206,0,254),(73,17,0,254),(8,17,0,254),(8,17,0,165),(8,17,138,165),(103,17,138,165),(103,80,138,165),(103,80,138,4),(103,222,138,4),(103,152,138,4),(34,152,138,4),(34,152,181,4),(34,152,181,21),(34,71,181,21),(0,0,0,197),(0,213,0,197),(48,213,0,197),(165,213,0,197),(0,0,15,0),(232,0,15,0),(184,0,15,0),(184,0,15,13),(184,0,15,242),(184,0,141,242),(184,148,141,242),(184,205,141,242),(184,240,141,242),(184,240,141,42),(184,240,141,222),(184,254,141,222),(184,144,141,222),(67,144,141,222),(67,144,141,129),(67,144,141,194),(0,0,115,0),(0,0,77,0),(0,0,77,101),(0,36,77,101),(102,36,77,101),(0,0,74,0),(0,201,0,0),(0,64,0,0),(0,90,0,0),(0,90,0,240),(0,90,30,240),(61,90,30,240),(18,90,30,240),(18,90,45,240),(18,90,45,85),(18,229,45,85),(18,229,86,85),(18,229,31,85),(18,229,31,249),(229,229,31,249),(229,229,31,7),(229,1,31,7),(229,214,31,7),(229,70,31,7),(182,70,31,7),(182,70,32,7),(182,177,32,7),(182,177,32,75),(182,177,145,75),(0,0,0,20),(0,15,0,20),(0,15,14,20),(0,15,14,12),(41,15,14,12),(41,15,14,172),(41,15,194,172),(41,93,194,172),(203,93,194,172),(203,93,103,172),(203,20,103,172),(203,20,103,16),(203,20,15,16),(203,20,201,16),(0,0,0,225),(0,77,0,225),(0,77,218,225),(0,31,218,225),(0,31,218,76),(0,197,218,76),(0,197,218,46),(88,197,218,46),(88,200,218,46),(0,0,27,0),(0,0,27,163),(116,0,27,163),(116,0,27,144),(116,197,27,144),(116,197,202,144),(60,197,202,144),(60,242,202,144),(60,242,202,206),(0,244,0,0),(0,44,0,0),(66,44,0,0),(66,44,0,169),(0,0,0,125),(118,0,0,125),(219,0,0,125),(219,0,42,125),(219,0,58,125),(219,0,58,11),(219,0,58,103),(219,0,199,103),(162,0,199,103),(162,0,244,103),(162,202,244,103),(0,0,0,48),(0,0,238,48),(0,85,238,48),(0,85,134,48),(0,85,134,117),(211,85,134,117),(211,85,136,117),(211,234,136,117),(31,234,136,117),(53,234,136,117),(53,118,136,117),(53,95,136,117),(53,95,118,117),(67,95,118,117),(67,95,118,4),(67,95,118,244),(67,95,29,244),(67,148,29,244),(37,148,29,244),(37,148,69,244),(246,148,69,244),(109,148,69,244),(242,148,69,244),(242,148,130,244),(242,206,130,244),(242,243,130,244),(242,217,130,244),(242,66,130,244),(242,13,130,244),(242,66,130,244),(156,66,130,244),(156,65,130,244),(73,0,0,0),(0,0,0,44),(152,0,0,44),(152,167,0,44),(152,167,0,218),(152,167,60,218),(152,15,60,218),(152,78,60,218),(152,78,60,218),(152,78,60,241),(152,78,60,168),(152,78,60,76),(0,165,0,0),(0,165,209,0),(0,173,209,0),(0,127,209,0),(0,127,209,179),(189,127,209,179),(0,0,26,0),(0,242,26,0),(212,242,26,0),(212,87,26,0),(0,0,236,0),(0,0,236,114),(0,0,86,114),(0,0,153,114),(0,0,153,169),(0,0,0,30),(0,166,0,30),(52,166,0,30),(52,166,78,30),(52,166,31,30),(42,166,31,30),(42,166,31,153),(42,166,234,153),(42,166,46,153),(42,166,46,6),(191,166,46,6),(151,166,46,6),(0,0,83,0),(0,41,0,0),(0,41,144,0),(0,41,144,127),(0,112,144,127),(0,116,144,127),(0,116,169,127),(78,0,0,0),(78,0,246,0),(78,0,246,164),(152,0,246,164),(152,114,246,164),(152,114,244,164),(152,114,131,164),(20,114,131,164),(20,114,238,164),(20,114,248,164),(20,114,248,252),(102,0,0,0),(39,0,0,0),(39,0,0,193),(39,211,0,193),(39,211,177,193),(92,211,177,193),(92,7,177,193),(92,7,177,46),(92,7,177,122),(92,7,177,92),(92,7,11,92),(92,204,11,92),(92,204,11,185),(58,204,11,185),(98,204,11,185),(98,204,31,185),(98,204,31,158),(126,0,0,0),(126,0,167,0),(105,0,167,0),(105,0,167,51),(105,0,191,51),(105,0,243,51),(105,85,243,51),(105,85,243,223),(105,85,243,71),(105,146,243,71),(105,73,243,71),(88,73,243,71),(88,73,161,71),(221,73,161,71),(0,0,23,0),(0,0,254,0),(0,0,254,101),(0,0,254,58),(0,0,254,48),(0,0,234,48),(0,0,113,48),(15,0,113,48),(15,160,113,48),(15,160,113,187),(15,160,95,187),(15,44,95,187),(210,44,95,187),(57,44,95,187),(57,44,80,187),(57,44,68,187),(57,44,83,187),(57,44,30,187),(57,44,163,187),(57,154,163,187),(0,102,0,0),(0,102,10,0),(0,102,10,147),(64,0,0,0),(64,0,141,0),(90,0,141,0),(90,0,141,152),(90,0,236,152),(90,0,74,152),(0,196,0,0),(0,196,0,242),(0,196,0,229),(225,0,0,0),(225,0,66,0),(225,0,31,0),(176,0,31,0),(35,0,0,0),(32,0,0,0),(32,0,203,0),(162,0,203,0),(0,0,245,0),(0,0,53,0),(213,0,53,0),(213,176,53,0),(213,176,53,28),(213,102,53,28),(213,102,53,209),(213,102,53,185),(213,102,53,113),(213,236,53,113),(213,236,53,125),(213,236,53,181),(0,236,53,181),(0,77,53,181),(0,77,87,181),(0,0,0,108),(0,127,0,108),(196,127,0,108),(196,127,0,140),(196,5,0,140),(186,5,0,140),(186,5,0,253),(186,5,44,253),(186,5,44,190),(186,5,107,190),(56,5,107,190),(56,5,107,216),(217,0,0,0),(217,223,0,0),(217,223,0,11),(217,223,200,11),(217,223,171,11),(94,223,171,11),(94,223,171,198),(94,30,171,198),(94,30,225,198),(204,30,225,198),(204,75,225,198),(204,75,225,49),(204,191,225,49),(165,0,0,0),(165,0,138,0),(226,0,138,0),(0,0,88,0),(0,0,205,0),(0,0,205,156),(0,0,233,156),(194,0,0,0),(194,0,182,0),(194,0,54,0),(210,0,54,0),(210,0,54,119),(210,0,54,43),(210,0,46,43),(17,0,46,43),(17,0,145,43),(17,0,145,166),(17,0,145,102),(17,29,145,102),(17,29,145,52),(17,29,7,52),(57,29,7,52),(138,29,7,52),(138,184,7,52),(70,184,7,52),(70,184,7,0),(70,180,7,0),(70,178,7,0),(0,0,100,0),(0,0,177,0),(0,0,177,45),(0,0,141,45),(176,0,141,45),(176,0,78,45),(176,166,78,45),(176,166,22,45),(176,166,22,106),(149,0,0,0),(105,0,0,0),(105,0,0,216),(105,0,92,216),(105,0,92,155),(92,0,92,155),(92,0,61,155),(92,0,169,155),(92,0,232,155),(84,0,232,155),(84,212,232,155),(84,122,232,155),(84,113,232,155),(84,113,232,57),(84,113,232,247),(84,113,232,244),(84,113,106,244),(84,113,238,244),(84,113,238,158),(0,0,0,169),(0,0,74,169),(0,253,74,169),(31,253,74,169),(31,225,74,169),(31,225,74,189),(46,225,74,189),(46,225,207,189),(46,99,207,189),(46,35,207,189),(46,5,207,189),(46,5,207,131),(46,175,207,131),(46,175,142,131),(74,175,142,131),(74,175,90,131),(74,14,90,131),(74,220,90,131),(59,220,90,131),(59,181,90,131),(59,181,90,105),(59,156,90,105),(59,156,53,105),(59,134,53,105),(59,134,53,21),(59,134,213,21),(236,134,213,21),(236,21,213,21),(24,21,213,21),(47,21,213,21),(47,21,213,247),(131,21,213,247),(131,21,213,25),(131,21,184,25),(131,21,26,25),(131,91,26,25),(131,88,26,25),(131,88,181,25),(131,88,181,12),(131,150,181,12),(131,150,15,12),(11,150,15,12),(11,150,15,123),(11,121,15,123),(11,121,15,156),(190,121,15,156),(190,121,194,156),(243,121,194,156),(243,121,44,156),(88,0,0,0),(88,0,38,0),(88,117,38,0),(88,117,32,0),(88,117,250,0),(88,117,250,96),(213,117,250,96),(213,243,250,96),(213,80,250,96),(0,106,0,0),(0,106,0,51),(0,106,0,36),(0,106,39,36),(58,0,0,0),(58,137,0,0),(58,64,0,0),(58,64,0,226),(58,64,136,226),(58,64,201,226),(58,24,201,226),(58,183,201,226),(210,183,201,226),(131,183,201,226),(60,183,201,226),(60,174,201,226),(60,96,201,226),(60,142,201,226),(151,142,201,226),(114,142,201,226),(114,142,237,226),(114,237,237,226),(114,237,135,226),(114,237,246,226),(114,237,31,226),(114,237,34,226),(114,237,34,29),(114,237,34,188),(114,237,43,188),(114,237,43,252),(114,237,184,252),(114,237,184,22),(88,237,184,22),(179,237,184,22),(0,0,0,29),(171,0,0,29),(171,26,0,29),(179,26,0,29),(179,105,0,29),(179,105,92,29),(179,105,155,29),(179,105,155,222),(179,155,155,222),(76,0,0,0),(219,0,0,0),(219,0,0,105),(219,14,0,105),(0,0,0,182),(0,56,0,182),(0,56,47,182),(0,225,47,182),(162,225,47,182),(162,225,168,182),(162,225,42,182),(162,225,89,182),(80,225,89,182),(0,5,0,0),(0,74,0,0),(0,74,51,0),(0,74,51,55),(0,74,71,55),(0,74,194,55),(188,0,0,0),(188,0,8,0),(0,0,147,0),(0,233,147,0),(0,233,147,125),(0,0,0,20),(48,0,0,0),(16,0,0,0),(16,147,0,0),(247,147,0,0),(0,0,191,0),(22,0,191,0),(22,168,191,0),(22,197,191,0),(22,197,191,192),(22,229,191,192),(188,0,0,0),(188,0,0,127),(101,0,0,127),(19,0,0,127),(19,0,84,127),(176,0,84,127),(176,36,84,127),(176,36,84,49),(176,36,84,140),(0,0,0,215),(0,0,31,215),(0,36,31,215),(0,36,31,100),(0,228,31,100),(0,228,192,100),(0,0,0,145),(120,0,0,0),(62,0,0,0),(62,0,0,131),(210,0,0,131),(210,174,0,131),(160,174,0,131),(160,174,2,131),(160,174,2,94),(73,174,2,94),(73,174,2,176),(113,174,2,176),(113,186,2,176),(31,186,2,176),(0,0,28,0),(52,0,28,0),(52,0,28,16),(0,165,0,0),(187,165,0,0),(187,165,0,37),(187,165,155,37),(187,165,44,37),(187,165,60,37),(187,165,108,37),(187,165,25,37),(216,165,25,37),(216,165,25,30),(216,98,25,30),(216,139,25,30),(0,0,0,6),(0,0,0,158),(92,0,0,158),(92,142,0,158),(219,0,0,0),(29,0,0,0),(170,0,0,0),(170,0,0,42),(170,0,149,42),(170,0,62,42),(170,0,148,42),(170,0,203,42),(170,75,203,42),(170,75,236,42),(170,75,236,228),(140,0,0,0),(118,0,0,0),(0,0,204,0),(98,0,204,0),(0,0,135,0),(0,0,135,171),(0,174,135,171),(247,174,135,171),(69,174,135,171),(93,0,0,0),(0,44,0,0),(0,182,0,0),(136,182,0,0),(136,210,0,0),(240,0,0,0),(151,0,0,0),(0,0,0,10),(0,0,66,10),(0,53,66,10),(39,0,0,0),(39,0,130,0),(39,0,70,0),(39,81,70,0),(39,81,70,20),(231,81,70,20),(231,81,196,20),(231,81,251,20),(231,81,149,20),(231,81,149,99),(231,81,176,99),(231,175,176,99),(231,175,176,111),(231,175,146,111),(231,96,146,111),(241,96,146,111),(61,96,146,111),(61,96,146,56),(163,96,146,56),(163,96,243,56),(153,96,243,56),(86,96,243,56),(86,96,243,165),(59,96,243,165),(59,96,243,35),(0,0,0,115),(0,113,0,115),(0,113,0,15),(226,113,0,15),(226,113,0,245),(226,113,0,179),(226,109,0,179),(226,109,0,167),(226,144,0,167),(226,144,159,167),(226,213,159,167),(226,213,172,167),(226,174,172,167),(226,57,172,167),(226,202,172,167),(0,0,0,233),(24,0,0,0),(24,56,0,0),(24,56,0,212),(24,226,0,212),(72,226,0,212),(72,226,0,38),(72,143,0,38),(72,143,0,41),(72,143,83,41),(72,143,83,229),(72,143,83,222),(72,143,99,222),(35,0,0,0),(35,129,0,0),(35,129,0,123),(35,129,0,254),(35,129,50,254),(35,129,50,233),(245,129,50,233),(245,129,23,233),(245,29,23,233),(241,29,23,233),(241,29,237,233),(241,29,237,142),(228,29,237,142),(0,227,0,0),(0,234,0,0),(109,0,0,0),(109,0,77,0),(109,0,77,175),(109,0,77,77),(109,0,77,10),(224,0,77,10),(184,0,77,10),(184,33,77,10),(184,33,164,10),(184,33,226,10),(0,0,61,0),(132,0,61,0),(132,0,43,0),(7,0,43,0),(7,82,43,0),(7,164,43,0),(7,88,43,0),(7,88,212,0),(138,88,212,0),(153,88,212,0),(153,88,124,0),(227,88,124,0),(16,88,124,0),(16,171,124,0),(16,171,124,24),(16,171,124,24),(225,171,124,24),(225,171,119,24),(225,171,119,207),(9,171,119,207),(114,0,0,0),(38,0,0,0),(240,0,0,0),(115,0,0,0),(115,82,0,0),(115,82,0,162),(115,82,224,162),(115,82,7,162),(115,82,235,162),(24,82,235,162),(61,82,235,162),(61,82,235,23),(112,82,235,23),(112,26,235,23),(112,106,235,23),(112,106,51,23),(112,106,238,23),(122,106,238,23),(137,106,238,23),(137,106,71,23),(137,60,71,23),(36,0,0,0),(36,0,175,0),(36,0,65,0),(36,170,65,0),(36,170,65,70),(36,170,65,215),(220,170,65,215),(220,170,65,137),(185,170,65,137),(185,170,65,33),(185,170,94,33),(185,170,94,217),(252,170,94,217),(252,170,94,85),(252,170,35,85),(252,170,35,37),(252,170,14,37),(252,170,43,37),(252,170,55,37),(105,170,55,37),(105,170,55,240),(105,170,7,240),(105,170,7,82),(105,169,7,82),(105,169,7,213),(34,169,7,213),(34,66,7,213),(34,66,7,40),(34,8,7,40),(34,8,7,27),(103,8,7,27),(103,133,7,27),(0,0,0,156),(0,0,0,152),(0,28,0,152),(0,28,0,116),(0,28,95,116),(0,28,6,116),(0,47,6,116),(0,47,76,116),(75,47,76,116),(75,142,76,116),(75,142,76,168),(88,142,76,168),(88,76,76,168),(88,76,76,206),(178,76,76,206),(178,212,76,206),(178,212,207,206),(178,212,207,178),(178,212,207,12),(178,151,207,12),(178,219,207,12),(178,12,207,12),(178,12,67,12),(178,12,67,18),(61,12,67,18),(61,12,67,38),(61,179,67,38),(61,179,67,73),(61,124,67,73),(61,223,67,73),(61,34,67,73),(202,34,67,73),(202,34,67,24),(202,52,67,24),(202,10,67,24),(202,10,13,24),(202,151,13,24),(202,173,13,24),(202,216,13,24),(202,216,13,105),(79,216,13,105),(79,190,13,105),(79,194,13,105),(79,194,118,105),(161,194,118,105),(246,194,118,105),(246,194,126,105),(246,194,164,105),(246,194,124,105),(42,194,124,105),(116,194,124,105),(116,194,124,4),(116,194,124,231),(116,194,124,126),(54,194,124,126),(54,194,27,126),(54,194,199,126),(232,194,199,126),(232,194,87,126),(232,62,87,126),(116,62,87,126),(222,0,0,0),(222,0,203,0),(218,0,203,0),(218,0,180,0),(218,145,180,0),(218,145,180,15),(218,145,119,15),(218,200,119,15),(191,200,119,15),(191,200,119,3),(191,167,119,3),(191,167,225,3),(191,139,225,3),(191,139,225,131),(63,139,225,131),(210,139,225,131),(210,151,225,131),(210,151,41,131),(83,151,41,131),(0,0,151,0),(0,0,183,0),(0,0,183,148),(0,0,183,122),(0,0,76,122),(168,0,76,122),(168,0,141,122),(0,0,129,0),(0,40,129,0),(230,40,129,0),(230,40,129,80),(167,40,129,80),(167,40,129,29),(126,40,129,29),(234,40,129,29),(234,46,129,29),(234,46,129,88),(234,46,129,138),(142,46,129,138),(142,46,169,138),(93,46,169,138),(93,200,169,138),(189,200,169,138),(189,200,169,94),(189,200,169,153),(189,139,169,153),(189,254,169,153),(189,254,169,240),(32,254,169,240),(32,254,169,180),(32,254,151,180),(32,254,199,180),(32,254,19,180),(32,45,19,180),(32,45,51,180),(32,45,51,8),(32,45,51,128),(32,45,93,128),(75,0,0,0),(166,0,0,0),(166,0,0,63),(0,149,0,0),(0,149,0,222),(0,149,0,21),(0,149,0,31),(0,149,0,47),(68,149,0,47),(68,149,138,47),(68,127,138,47),(0,171,0,0),(0,171,0,80),(0,171,239,80),(0,18,239,80),(0,18,67,80),(0,18,67,73),(0,18,67,231),(0,18,96,231),(0,18,96,72)
	);

	SIGNAL do_reset : std_logic_vector(0 TO N_EVENTS - 1) := "1000000000000000001100000000000000100100100000000000010000000000000000000000000000000010000100000000100000000000010010000000000001001000000000000000000100000100000000000001000000000000001000100010100000000000000000000010000000000000000000000000100000000000000000101000000000000000000100001000000000000000000000010001000000000110000000000000000010110000100000000000000000000000000000100000000100000001000000000000000001000000100000000000000000000001000000000000000000000000000001000001000000101000000000000000001000000000001001000000000000000000000000000001000100000100000000000101000000101000000001000000000001000011010000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000001000000000100001000000001000000100010000010000010000000000000001011000000000001000001000000000000000000000000000000001000000000000000000000000000000000000000000000000100000000001000000000000000100000000000110000000100000100000000000100000000001100000100100001000100000000000000000000010010000010000000100000000000000000000000000010000000000000001000000000000000000000001000000000000000000000000000011000000010000010000000100000010000000010000000000000011100000000000000100001000110001000000000000000000000000000010000000000000000000000000000100100000000000001000000000100000000010000000000000100000000000000000000000000000000000000000000000000001000100000000000000000000001000001000000000000000000010000000000000000000000000100001000000000000000000000000000000000000000000000000000010000000000010000000000000000010001000000000000000000010000100000000000000000000000000010100000000000100000001001000000000000000001000000000000001000000000000100000000000000000000000000000010010000000000000000000000100000010000000000000100000000000000000000000000000000000000001000000000000000000010100001000000000000000000110000000000000000000000000000110010000000000110000000000000000000000000000001000000100000000000000000000000100000000000010000010101000000000000100000100000011000101000000000000000000000000000000000000000000001000000100000000000000000100000000000000000000000000000110000100000000100001000000000010000010000000000000000000000000000000000000000100000000001010000100000000000000000000001000000000000000000000000000100000000000000000100000000000100000010000000000000000000000000000000000000001000000000000000000000010010000000000000000000000000000000000000000000100000110000000000001000000000000000100000001010001000000000000000000100000000000000000000000000000000100010000000000000000000000000000100000000000000000000000000000110000000000000001110000000000000000000010000000100000000000000000000100010000000100010000000000000000000000000000000000000000000000000001010100010000010000000000000000011000000000000000000000001010000000100000000000000000100001000000000000000000000000010000000000000000000000000000000001000000000100000000010000000100000000000100001000000000000000000000000000000000000001000000100100000101000000000000000000000010000100010000000000001000000100000010000000000100000010010000110000000000000000000000000000000000000100000000000000000000000000000001000000001000100000000000000000000000000000000000001000000000000000000000100000000000000000000000000000010000010001000010000000000000000011000000010000000000000000000001000000010000000000001000000000000100000000000000100000000000000000000000000000000000000000000000000000010000000000001000000000000000001000000000000000000100000000011000000000000000000000000000100010000000000100000000000000000000000001001100000100001000000100000000000001010000100010100010000000000000010000000000000000000110000000000000000000000000000000100000000010001000001010000000000000000001000000000001000000000000000000000000100000000000000000000000001010000000000100010010000000000000000000000000000000000001000000000000100001000001100000001000000000000000000000000100010000000100000010000000000000000001000000001000000000000000000001000000100000000000000000000000001000001000100010000010000000000000000000000000000000000010000000000001000000000100000000000000000000000000000000001000000000000000100000100010000010000110000000000100001000000000000000000100010000000000001000000000000000000010000000000000000000000000100010000000000001000000000000000000000100000000010000000000000000000000000000000010000000000000000001000000000001010000001000000000000000010010000001000000010000000010000000000000000000000010000000000000000000010000000001000000000000000000000100000010001000000101000000000101000000010000000000000000000000000000000000011000100010110000000000100000000000001000100000000101000000000000000000010000000000000100001000011000000000001000010000000000000000010000000000000000000000000000000101000000000000000001000000000001000000000000000000000000000000001000000001010000000000000001100000001000010010000000000000100000100000000100010100011000000000000000000000000000000000000000000000000000000000010000000000000000000100000000000000000000100000100000000000000000000010000101011000000000000000000000000000000000000001100000000001100000000000000010010000000000000000000100100000000100010000000001010000000000000000001010000000000100000010000000000000000001100100100001100000000000000000010000000000000000000001000000000000010000000000000000000001000000000000000010001000010000000000100000000000001000000100000000100000000000000000000000000000001000000000010010000001000000000010000001000000011101000000000000000000000000000100000010001000000000000010000000001000000000000010000000000010001000000000000010000010000000100000010000101000010000000000000000000000000000010000000000101000000000000100000000000010001000001000000100000000100000000000000000000010000000000000000000000000000000001001000000000000100000000000001000000000001101000000000000000000000100100000000000000000000010000000010000000000000010100000001000100100000000000000001000000000010000010000010000000000000000010010000000000000000000100000000100000000100000000000000000000001000000000010000000000000000001000000001010000001010000000000000001010000000001010000000000000000000000000001000000000000001000000000000000000000010010000000000000010000000001000000100000000000000000000010000000000000001000100000000100000000000001010000101000000000000000000000000000000000010000000100000000000000000100000001000000000000000000000010000000010000000000010000000000100001001000000100000000010000010000000000000000100000000000000000000000000000010000000000100010000000000000000100000100000000000100000000110001010000000000000100000010000000001010010000000000000100000000010001000000000010000000010000000000000000000000100001010000000000000100000000001010000000000000000000000000001000000000000000000000000000001000001000010000000000100000000000000000000000000000000000000100000000010001000000000100000100000100000000000000000000000000000000101100000000000000000000001001000000000000000000000000000000000000000000000001000000000110001000101000000000000000100000100000000000100010000000000000101000000000001000000000000000100000000000101000000000000000000000100010000001000000110000000000000100000000000010000000000000001000000000010000000000101000001000000000000000100000000000000000001000000000000000000000000001000000000000000000000000010000000000000000000000000000000000000000000000010100000010001000000000000000000000110000001001000000000000100000000000000000000000001010000100000000000000000000000000000010000000000000000000000000000010000000000000000000010000000000000000001000000100010010000000001000000000001000000000000000000010000000000000000000000010000000100000000000000100000000100000010000010000000000100111001000000010000010000010000100000000000000000000000000000001000100000010000000010100010000000000001000000001000000000000000010000000010000000000000000001001000000000000000000000100000000100000000000000010000000100001000000100000000101000000010000110010000010000000000000000011000100000000000000000000000000000000000000010000000000000000000000100000010100000000000100000001000000000000000000000000000000100000000000000000000001010000110000000000000000000000000000000000000000000000000000000000001010000101000000001100001000000000000010000000000000000000000000010000000101000000000000010001000100100000010000000000001000001000000101000000000000000000000000000000000000000000000100000000000000100000000000000000000000000000100000000001010000000000000000000000000000000010001000010000010011000000000000000000000000010000000000001000000010001000100000010100100110100000000100000000101000000100100000000100001000000001000000000000010000100000000000100000000000000100000000100000000000000000000000000000000000000000000000000000000000000000000011100000000000100000000000000001000000000000010000000000000000100000000000000001000000001010000010000001000000000001000000000000100000000010000000000000000000000000000000001000000000010001100000000000000000000101000000000010001000000110000000000000000000000000000000000000010100000000000001000000000000000000000000000001000100100010000000000000100000000000000010000010000000100100000000000000000001000010000000000000000000000000000000000000001000000000000000010000000000000000010000000000000001000000000000000101000000000100000000101010001000000000000000000100010000000000000001000011000000000000000000000010000000000000100000000100000000100010000000000100000000000000000000000000000001100000000001000001000100001000000000001100000100000000001000000000000000010000000000000100000000000000000001001000001001000100010000000000000010000000000010000000000001001000100000000000000000000100000000100000000000000000010000000000000000000000000000000000000000000000001000000001000100000000000000000000000000000100000000100010000000010000010100110001000001000000001000001100000000000010010000000000010001000000000010101000011000101001000000000000000000000000100000000000000110000000000010000000000001010000000001000000000000000000010000000000000000000010000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000010000000000000000001000000100000000000000000000000000000010010000000100000000";

	TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL RAM : ram_type := (
		11 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		15 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		16 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		25 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		27 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		28 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		40 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		52 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		59 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		60 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		65 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		71 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		74 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		81 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		83 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		101 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		102 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		120 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		125 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		139 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		146 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		154 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		158 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		161 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		162 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		167 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		168 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		187 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		192 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		204 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		208 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		211 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		220 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		223 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		225 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		245 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		250 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		252 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		255 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		256 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		259 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		267 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		289 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		290 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		299 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		314 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		318 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		325 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		344 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		351 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		354 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		359 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		371 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		378 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		380 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		382 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		387 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		400 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		405 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		408 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		410 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		427 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		428 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		440 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		452 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		456 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		457 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		461 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		464 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		466 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		482 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		491 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		506 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		512 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		513 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		516 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		519 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		526 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		532 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		542 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		547 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		550 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		557 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		560 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		562 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		565 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		567 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		571 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		582 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		590 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		604 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		611 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		622 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		638 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		651 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		652 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		674 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		678 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		679 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		690 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		692 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		698 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		699 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		701 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		705 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		708 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		729 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		739 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		741 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		745 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		746 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		761 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		775 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		779 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		780 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		791 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		799 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		802 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		813 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		819 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		820 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		844 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		855 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		856 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		858 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		862 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		867 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		873 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		874 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		878 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		879 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		902 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		903 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		906 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		912 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		917 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		926 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		933 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		936 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		943 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		951 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		955 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		960 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		970 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		989 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		993 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		997 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		1014 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		1015 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		1030 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		1035 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		1060 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		1065 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		1066 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		1074 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		1083 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		1094 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		1101 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		1107 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		1112 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		1127 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		1139 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		1140 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		1154 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		1156 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		1163 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		1173 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		1174 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		1176 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		1181 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		1204 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		1226 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		1230 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		1241 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		1246 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		1251 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		1262 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		1274 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		1282 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		1305 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		1310 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		1312 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		1316 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		1326 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		1333 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		1348 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		1357 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		1373 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		1387 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		1394 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		1410 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		1415 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		1426 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		1430 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		1434 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		1455 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		1456 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		1459 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		1461 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		1462 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		1490 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		1491 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		1498 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		1507 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		1508 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		1512 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		1517 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		1519 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		1536 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		1537 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		1545 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		1546 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		1547 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		1552 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		1557 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		1561 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		1572 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		1574 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		1587 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		1588 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		1593 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		1598 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		1604 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		1616 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		1626 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		1638 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		1639 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		1642 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		1646 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		1652 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		1656 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		1661 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		1663 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		1666 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		1681 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		1682 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		1683 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		1690 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		1700 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		1715 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		1717 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		1727 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		1732 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		1745 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		1751 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		1753 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		1782 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		1793 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		1795 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		1805 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		1807 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		1814 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		1819 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		1830 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		1831 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		1843 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		1844 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		1845 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		1848 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		1849 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		1850 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		1859 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		1865 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		1878 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		1880 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		1881 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		1904 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		1907 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		1916 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		1918 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		1923 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		1929 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		1935 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		1949 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		1953 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		1977 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		1979 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		1986 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		1997 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		1999 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		2007 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		2013 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		2019 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		2023 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		2027 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		2030 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		2039 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		2041 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		2052 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		2074 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		2075 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		2078 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		2079 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		2080 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		2083 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		2090 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		2139 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		2140 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		2144 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		2149 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		2164 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		2167 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		2171 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		2175 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		2188 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		2189 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		2195 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		2198 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		2202 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		2226 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		2229 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		2231 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		2242 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		2256 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		2267 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		2279 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		2298 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		2308 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		2310 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		2320 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		2331 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		2364 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		2373 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		2379 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		2397 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		2408 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		2433 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		2444 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		2457 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		2461 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		2471 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		2473 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		2487 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		2490 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		2495 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		2498 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		2505 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		2524 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		2528 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		2540 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		2546 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		2551 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		2555 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		2575 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		2577 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		2582 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		2585 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		2586 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		2588 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		2598 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		2610 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		2620 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		2621 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		2628 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		2636 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		2646 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		2652 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		2665 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		2693 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		2710 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		2717 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		2726 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		2732 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		2738 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		2756 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		2759 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		2760 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		2765 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		2769 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		2770 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		2776 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		2778 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		2783 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		2785 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		2786 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		2804 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		2809 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		2813 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		2821 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		2824 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		2825 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		2832 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		2844 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		2863 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		2870 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		2873 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		2875 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		2880 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		2907 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		2911 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		2913 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		2922 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		2923 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		2928 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		2935 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		2936 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		2940 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		2942 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		2966 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		2968 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		2973 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		2977 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		2989 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		3004 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		3007 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		3008 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		3011 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		3020 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		3031 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		3039 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		3043 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		3058 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		3067 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		3072 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		3080 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		3107 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		3108 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		3123 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		3132 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		3133 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		3134 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		3135 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		3140 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		3156 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		3160 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		3169 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		3171 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		3177 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		3178 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		3181 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		3197 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		3199 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		3200 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		3203 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		3212 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		3214 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		3229 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		3234 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		3236 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		3253 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		3254 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		3260 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		3268 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		3274 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		3275 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		3276 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		3281 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		3286 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		3288 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		3308 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		3316 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		3322 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		3335 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		3336 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		3338 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		3340 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		3341 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		3347 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		3350 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		3352 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		3393 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		3405 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		3407 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		3408 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		3420 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		3423 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		3427 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		3436 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		3439 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		3440 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		3454 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		3459 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		3465 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		3475 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		3481 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		3490 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		3491 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		3516 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		3523 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		3540 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		3542 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		3567 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		3573 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		3575 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		3578 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		3585 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		3590 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		3596 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		3599 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		3603 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		3613 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		3617 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		3623 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		3632 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		3633 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		3638 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		3642 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		3646 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		3649 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		3650 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		3652 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		3654 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		3661 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		3663 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		3670 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		3677 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		3678 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		3683 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		3694 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		3699 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		3708 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		3713 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		3729 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		3733 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		3743 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		3755 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		3756 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		3760 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		3773 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		3775 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		3788 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		3790 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		3797 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		3800 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		3801 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		3803 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		3814 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		3815 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		3821 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		3835 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		3838 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		3846 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		3847 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		3852 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		3858 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		3861 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		3876 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		3877 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		3888 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		3897 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		3906 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		3907 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		3909 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		3910 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		3911 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		3912 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		3917 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		3926 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		3930 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		3932 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		3934 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		3951 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		3953 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		3956 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		3965 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		3972 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		3973 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		3985 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		3992 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		3997 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		4002 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		4003 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		4005 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		4012 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		4022 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		4025 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		4026 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		4036 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		4037 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		4049 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		4053 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		4054 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		4057 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		4059 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		4072 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		4077 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		4087 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		4088 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		4089 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		4096 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		4106 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		4108 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		4120 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		4121 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		4130 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		4138 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		4143 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		4145 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		4152 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		4156 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		4160 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		4162 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		4172 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		4175 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		4176 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		4178 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		4195 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		4204 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		4206 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		4207 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		4219 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		4220 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		4226 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		4232 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		4235 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		4242 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		4248 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		4272 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		4278 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		4289 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		4296 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		4309 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		4312 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		4313 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		4316 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		4324 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		4330 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		4331 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		4333 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		4336 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		4345 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		4378 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		4391 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		4398 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		4405 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		4407 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		4416 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		4417 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		4425 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		4430 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		4434 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		4489 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		4494 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		4495 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		4498 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		4500 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		4501 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		4502 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		4533 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		4537 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		4544 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		4547 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		4551 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		4563 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		4566 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		4579 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		4580 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		4581 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		4582 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		4583 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		4584 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		4585 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		4587 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		4595 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		4612 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		4615 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		4616 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		4639 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		4649 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		4670 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		4682 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		4683 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		4697 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		4720 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		4737 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		4742 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		4743 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		4749 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		4750 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		4753 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		4759 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		4761 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		4763 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		4769 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		4770 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		4771 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		4775 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		4777 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		4781 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		4784 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		4785 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		4791 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		4799 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		4800 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		4852 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		4862 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		4871 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		4874 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		4876 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		4887 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		4889 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		4894 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		4909 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		4914 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		4916 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		4930 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		4938 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		4944 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		4945 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		4948 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		4949 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		4957 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		4965 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		4966 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		4972 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		4977 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		4986 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		4989 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		4997 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		5003 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		5009 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		5022 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		5031 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		5035 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		5040 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		5063 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		5067 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		5068 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		5074 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		5119 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		5122 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		5131 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		5143 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		5166 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		5169 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		5186 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		5187 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		5195 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		5209 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		5232 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		5235 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		5239 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		5248 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		5254 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		5260 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		5270 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		5273 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		5274 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		5277 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		5278 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		5284 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		5290 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		5291 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		5305 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		5308 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		5315 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		5320 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		5328 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		5330 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		5337 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		5343 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		5348 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		5350 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		5362 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		5373 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		5376 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		5380 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		5389 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		5396 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		5401 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		5407 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		5408 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		5413 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		5421 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		5427 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		5430 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		5431 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		5445 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		5448 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		5449 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		5457 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		5472 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		5475 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		5480 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		5489 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		5501 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		5510 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		5536 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		5537 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		5545 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		5552 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		5563 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		5564 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		5577 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		5579 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		5591 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		5593 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		5597 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		5603 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		5605 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		5612 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		5615 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		5617 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		5623 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		5638 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		5640 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		5647 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		5671 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		5674 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		5682 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		5718 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		5720 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		5721 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		5722 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		5724 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		5731 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		5732 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		5734 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		5744 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		5748 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		5750 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		5760 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		5762 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		5769 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		5772 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		5776 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		5778 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		5786 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		5805 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		5808 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		5813 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		5818 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		5819 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		5830 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		5839 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		5843 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		5868 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		5875 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		5877 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		5880 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		5888 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		5899 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		5901 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		5910 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		5916 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		5919 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		5921 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		5927 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		5934 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		5938 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		5945 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		5946 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		5948 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		5949 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		5952 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		5954 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		5963 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		5979 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		5995 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		5996 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		6008 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		6027 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		6042 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		6053 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		6054 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		6060 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		6063 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		6066 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		6072 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		6079 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		6088 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		6092 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		6093 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		6096 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		6106 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		6119 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		6131 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		6141 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		6144 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		6158 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		6159 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		6171 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		6172 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		6180 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		6192 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		6204 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		6207 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		6216 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		6218 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		6246 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		6259 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		6261 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		6267 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		6269 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		6272 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		6296 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		6297 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		6299 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		6306 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		6313 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		6317 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		6326 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		6336 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		6338 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		6347 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		6360 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		6362 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		6363 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		6365 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		6369 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		6370 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		6387 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		6388 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		6396 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		6403 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		6413 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		6422 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		6435 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		6437 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		6447 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		6477 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		6482 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		6484 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		6485 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		6491 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		6499 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		6506 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		6512 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		6517 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		6530 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		6531 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		6533 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		6546 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		6554 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		6560 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		6577 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		6584 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		6587 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		6590 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		6604 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		6622 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		6624 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		6634 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		6635 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		6642 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		6660 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		6663 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		6664 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		6678 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		6684 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		6685 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		6687 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		6701 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		6714 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		6722 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		6728 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		6765 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		6766 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		6772 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		6778 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		6787 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		6796 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		6803 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		6813 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		6815 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		6816 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		6818 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		6823 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		6866 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		6870 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		6876 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		6886 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		6899 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		6906 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		6907 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		6916 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		6919 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		6921 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		6923 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		6927 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		6950 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		6952 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		6972 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		6987 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		6991 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		7001 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		7004 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		7010 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		7018 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		7019 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		7021 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		7046 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		7047 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		7049 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		7052 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		7076 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		7078 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		7087 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		7105 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		7106 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		7107 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		7124 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		7132 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		7133 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		7140 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		7143 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		7145 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		7146 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		7147 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		7149 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		7150 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		7158 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		7161 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		7176 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		7179 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		7181 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		7184 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		7185 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		7213 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		7216 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		7220 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		7228 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		7243 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		7247 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		7252 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		7254 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		7261 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		7268 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		7270 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		7281 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		7282 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		7286 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		7313 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		7316 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		7320 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		7346 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		7364 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		7373 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		7377 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		7397 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		7408 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		7413 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		7417 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		7423 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		7426 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		7437 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		7439 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		7463 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		7464 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		7467 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		7472 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		7475 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		7489 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		7492 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		7501 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		7502 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		7503 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		7513 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		7516 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		7522 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		7526 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		7527 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		7529 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		7535 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		7547 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		7549 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		7555 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		7559 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		7565 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		7569 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		7576 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		7583 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		7596 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		7598 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		7603 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		7608 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		7617 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		7652 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		7661 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		7665 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		7670 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		7676 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		7687 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		7694 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		7695 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		7718 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		7723 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		7733 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		7737 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		7741 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		7749 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		7756 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		7764 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		7775 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		7786 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		7791 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		7793 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		7795 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		7796 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		7805 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		7822 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		7825 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		7828 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		7829 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		7849 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		7852 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		7853 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		7860 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		7863 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		7864 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		7875 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		7877 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		7878 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		7893 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		7896 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		7901 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		7919 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		7921 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		7928 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		7936 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		7958 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		7959 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		7962 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		7970 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		7980 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		7984 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		7985 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		7991 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		8002 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		8006 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		8016 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		8032 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		8034 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		8048 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		8051 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		8060 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		8063 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		8065 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		8084 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		8085 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		8086 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		8097 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		8101 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		8102 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		8115 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		8126 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		8129 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		8136 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		8139 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		8144 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		8145 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		8146 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		8148 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		8151 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		8155 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		8163 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		8166 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		8174 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		8182 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		8183 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		8187 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		8194 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		8200 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		8205 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		8206 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		8213 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		8218 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		8232 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		8233 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		8240 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		8246 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		8247 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		8253 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		8262 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		8264 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		8292 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		8298 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		8299 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		8302 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		8303 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		8307 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		8309 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		8316 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		8325 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		8327 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		8328 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		8329 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		8333 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		8339 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		8344 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		8345 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		8355 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		8357 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		8359 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		8361 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		8362 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		8373 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		8386 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		8395 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		8405 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		8420 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		8429 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		8432 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		8434 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		8450 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		8457 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		8458 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		8459 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		8461 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		8462 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		8465 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		8470 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		8477 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		8489 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		8494 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		8496 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		8501 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		8510 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		8523 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		8531 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		8533 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		8546 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		8548 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		8555 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		8569 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		8581 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		8585 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		8594 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		8597 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		8598 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		8605 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		8607 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		8615 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		8616 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		8618 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		8624 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		8628 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		8641 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		8642 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		8643 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		8676 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		8682 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		8694 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		8697 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		8698 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		8704 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		8705 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		8712 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		8715 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		8723 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		8740 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		8741 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		8743 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		8770 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		8783 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		8790 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		8792 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		8816 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		8823 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		8830 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		8832 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		8841 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		8851 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		8855 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		8861 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		8863 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		8869 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		8876 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		8896 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		8900 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		8910 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		8926 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		8927 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		8960 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		8967 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		8968 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		8969 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		8983 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		8984 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		8995 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		9003 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		9010 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		9019 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		9020 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		9033 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		9053 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		9070 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		9083 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		9085 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		9094 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		9097 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		9098 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		9099 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		9103 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		9111 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		9116 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		9125 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		9138 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		9146 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		9152 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		9155 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		9170 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		9173 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		9181 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		9189 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		9192 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		9197 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		9198 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		9209 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		9212 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		9217 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		9229 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		9233 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		9235 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		9241 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		9242 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		9247 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		9255 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		9261 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		9265 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		9266 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		9282 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		9284 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		9287 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		9302 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		9306 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		9311 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		9318 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		9325 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		9327 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		9330 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		9332 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		9333 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		9339 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		9345 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		9358 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		9368 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		9382 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		9401 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		9408 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		9412 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		9415 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		9442 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		9445 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		9446 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		9450 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		9452 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		9457 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		9460 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		9470 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		9471 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		9473 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		9483 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		9486 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		9495 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		9497 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		9499 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		9502 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		9539 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		9554 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		9559 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		9560 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		9562 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		9575 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		9579 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		9580 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		9593 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		9598 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		9602 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		9603 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		9608 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		9609 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		9614 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		9617 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		9619 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		9620 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		9625 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		9631 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		9638 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		9641 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		9666 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		9678 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		9679 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		9681 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		9682 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		9712 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		9717 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		9721 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		9726 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		9727 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		9728 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		9731 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		9737 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		9741 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		9743 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		9752 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		9753 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		9756 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		9763 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		9770 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		9772 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		9774 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		9775 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		9779 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		9780 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		9786 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		9803 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		9811 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		9817 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		9818 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		9821 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		9826 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		9829 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		9830 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		9832 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		9840 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		9845 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		9849 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		9854 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		9860 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		9869 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		9874 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		9877 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		9879 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		9898 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		9901 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		9908 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		9916 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		9918 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		9922 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		9925 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		9931 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		9937 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		9949 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		9953 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		9956 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		9959 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		9963 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		9964 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		9967 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		9979 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		9983 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		9984 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		9986 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		9987 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		9992 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		9999 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		10003 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		10008 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		10012 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		10016 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		10020 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		10021 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		10022 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		10025 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		10026 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		10039 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		10045 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		10053 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		10054 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		10058 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		10075 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		10078 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		10080 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		10082 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		10085 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		10086 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		10090 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		10104 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		10108 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		10113 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		10122 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		10134 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		10135 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		10140 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		10147 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		10154 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		10159 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		10171 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		10181 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		10182 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		10185 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		10194 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		10195 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		10204 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		10206 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		10218 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		10232 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		10238 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		10243 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		10256 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		10259 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		10262 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		10264 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		10265 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		10266 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		10269 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		10275 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		10281 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		10284 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		10285 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		10287 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		10292 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		10302 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		10315 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		10321 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		10324 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		10329 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		10334 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		10336 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		10344 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		10352 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		10357 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		10362 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		10364 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		10377 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		10397 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		10402 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		10405 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		10409 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		10413 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		10415 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		10437 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		10440 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		10445 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		10460 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		10464 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		10465 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		10479 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		10487 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		10520 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		10522 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		10526 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		10529 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		10540 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		10541 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		10547 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		10561 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		10565 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		10566 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		10567 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		10571 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		10580 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		10584 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		10630 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		10631 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		10662 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		10666 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		10670 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		10673 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		10698 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		10703 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		10713 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		10726 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		10739 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		10743 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		10749 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		10755 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		10764 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		10778 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		10781 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		10797 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		10807 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		10808 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		10810 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		10814 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		10828 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		10833 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		10836 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		10846 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		10852 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		10855 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		10863 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		10873 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		10883 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		10898 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		10901 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		10902 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		10914 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		10918 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		10919 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		10925 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		10928 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		10930 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		10947 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		10959 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		10961 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		10965 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		10974 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		10975 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		10979 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		10990 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		10993 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		10997 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		11000 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		11001 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		11004 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		11014 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		11016 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		11019 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		11022 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		11028 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		11032 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		11037 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		11043 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		11053 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		11065 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		11067 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		11070 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		11075 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		11078 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		11087 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		11108 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		11109 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		11154 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		11159 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		11161 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		11163 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		11170 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		11173 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		11175 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		11181 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		11185 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		11186 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		11189 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		11191 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		11207 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		11212 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		11213 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		11226 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		11233 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		11254 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		11260 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		11261 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		11262 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		11271 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		11293 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		11301 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		11308 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		11313 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		11319 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		11323 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		11339 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		11363 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		11368 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		11369 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		11380 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		11398 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		11403 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		11410 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		11412 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		11422 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		11425 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		11430 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		11432 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		11435 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		11449 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		11452 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		11454 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		11461 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		11462 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		11468 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		11470 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		11471 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		11473 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		11479 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		11487 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		11512 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		11518 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		11526 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		11531 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		11532 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		11537 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		11544 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		11545 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		11561 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		11562 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		11566 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		11574 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		11585 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		11596 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		11602 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		11623 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		11625 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		11632 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		11646 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		11654 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		11656 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		11661 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		11669 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		11670 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		11671 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		11683 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		11685 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		11708 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		11714 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		11738 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		11745 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		11748 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		11779 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		11781 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		11800 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		11826 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		11834 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		11836 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		11837 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		11841 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		11843 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		11853 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		11861 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		11875 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		11876 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		11881 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		11902 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		11908 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		11914 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		11915 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		11917 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		11921 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		11933 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		11936 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		11937 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		11959 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		11962 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		11963 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		11968 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		11976 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		11979 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		11981 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		11985 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		11987 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		11988 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		11989 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		11991 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		11993 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		12000 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		12004 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		12021 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		12031 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		12037 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		12040 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		12051 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		12074 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		12080 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		12081 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		12093 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		12094 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		12097 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		12109 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		12111 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		12114 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		12118 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		12122 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		12125 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		12127 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		12134 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		12138 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		12139 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		12141 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		12147 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		12167 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		12173 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		12177 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		12185 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		12187 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		12188 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		12192 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		12197 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		12217 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		12226 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		12232 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		12256 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		12265 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		12268 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		12289 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		12292 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		12299 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		12300 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		12303 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		12328 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		12347 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		12348 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		12351 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		12360 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		12363 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		12376 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		12378 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		12394 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		12405 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		12406 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		12407 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		12412 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		12419 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		12422 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		12443 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		12447 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		12458 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		12464 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		12470 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		12488 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		12490 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		12497 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		12514 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		12515 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		12516 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		12526 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		12551 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		12556 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		12561 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		12563 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		12565 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		12567 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		12573 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		12575 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		12577 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		12586 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		12599 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		12605 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		12606 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		12610 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		12615 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		12626 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		12657 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		12662 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		12664 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		12666 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		12680 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		12681 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		12686 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		12700 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		12717 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		12719 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		12721 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		12731 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		12733 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		12737 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		12738 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		12744 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		12747 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		12748 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		12750 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		12756 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		12766 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		12775 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		12784 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		12785 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		12793 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		12798 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		12803 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		12804 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		12815 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		12816 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		12825 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		12826 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		12827 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		12828 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		12848 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		12864 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		12867 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		12880 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		12882 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		12885 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		12886 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		12890 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		12891 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		12917 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		12928 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		12930 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		12931 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		12937 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		12938 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		12954 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		12982 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		13001 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		13004 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		13007 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		13015 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		13019 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		13021 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		13023 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		13031 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		13033 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		13043 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		13045 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		13058 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		13059 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		13065 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		13066 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		13067 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		13080 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		13088 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		13089 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		13093 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		13101 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		13108 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		13109 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		13110 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		13126 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		13127 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		13134 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		13137 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		13138 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		13146 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		13147 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		13156 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		13159 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		13163 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		13183 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		13197 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		13218 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		13221 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		13222 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		13225 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		13228 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		13240 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		13247 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		13265 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		13269 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		13275 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		13277 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		13289 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		13313 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		13317 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		13337 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		13350 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		13351 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		13369 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		13372 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		13375 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		13391 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		13395 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		13411 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		13418 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		13426 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		13427 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		13434 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		13444 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		13447 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		13452 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		13458 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		13462 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		13469 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		13472 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		13477 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		13485 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		13487 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		13499 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		13501 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		13503 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		13508 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		13511 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		13518 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		13519 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		13525 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		13535 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		13546 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		13550 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		13554 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		13569 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		13575 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		13582 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		13592 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		13596 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		13604 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		13607 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		13613 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		13614 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		13625 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		13628 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		13639 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		13642 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		13657 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		13663 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		13665 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		13670 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		13676 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		13678 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		13685 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		13688 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		13694 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		13708 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		13710 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		13725 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		13727 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		13731 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		13737 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		13745 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		13748 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		13755 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		13760 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		13762 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		13771 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		13775 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		13781 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		13798 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		13801 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		13805 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		13807 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		13808 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		13824 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		13839 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		13841 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		13847 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		13848 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		13858 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		13862 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		13866 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		13868 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		13870 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		13876 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		13881 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		13885 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		13888 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		13889 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		13893 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		13901 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		13902 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		13912 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		13917 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		13918 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		13921 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		13926 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		13937 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		13941 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		13947 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		13970 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		13971 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		13990 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		14008 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		14018 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		14020 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		14025 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		14030 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		14036 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		14045 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		14052 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		14054 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		14055 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		14059 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		14066 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		14082 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		14085 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		14099 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		14109 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		14119 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		14139 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		14144 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		14145 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		14146 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		14172 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		14177 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		14180 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		14183 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		14187 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		14206 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		14207 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		14214 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		14240 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		14253 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		14260 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		14270 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		14272 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		14276 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		14278 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		14281 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		14282 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		14283 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		14300 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		14305 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		14307 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		14309 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		14349 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		14363 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		14365 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		14392 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		14393 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		14396 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		14403 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		14413 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		14417 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		14418 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		14425 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		14441 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		14443 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		14445 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		14454 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		14465 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		14471 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		14476 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		14480 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		14485 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		14490 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		14493 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		14498 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		14501 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		14514 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		14522 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		14526 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		14528 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		14533 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		14544 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		14545 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		14551 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		14552 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		14575 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		14579 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		14589 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		14595 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		14600 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		14602 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		14609 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		14619 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		14636 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		14642 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		14651 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		14653 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		14663 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		14679 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		14686 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		14711 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		14722 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		14727 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		14731 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		14734 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		14737 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		14742 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		14744 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		14770 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		14773 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		14778 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		14780 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		14781 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		14786 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		14787 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		14796 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		14803 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		14804 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		14810 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		14813 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		14817 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		14819 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		14824 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		14828 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		14840 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		14842 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		14843 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		14852 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		14855 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		14857 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		14861 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		14862 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		14864 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		14867 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		14870 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		14871 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		14882 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		14889 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		14894 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		14902 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		14912 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		14919 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		14920 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		14925 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		14940 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		14944 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		14949 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		14953 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		14957 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		14972 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		14983 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		15013 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		15019 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		15026 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		15029 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		15030 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		15033 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		15034 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		15036 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		15052 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		15059 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		15075 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		15087 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		15091 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		15093 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		15108 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		15111 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		15112 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		15113 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		15114 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		15116 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		15119 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		15131 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		15137 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		15142 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		15143 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		15154 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		15161 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		15171 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		15187 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		15189 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		15215 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		15228 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		15229 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		15233 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		15237 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		15247 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		15250 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		15258 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		15263 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		15267 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		15275 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		15278 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		15281 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		15282 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		15287 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		15292 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		15294 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		15318 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		15321 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		15325 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		15337 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		15338 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		15340 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		15350 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		15364 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		15388 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		15390 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		15393 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		15398 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		15399 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		15403 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		15414 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		15420 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		15421 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		15424 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		15433 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		15444 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		15457 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		15463 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		15472 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		15473 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		15490 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		15518 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		15526 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		15534 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		15535 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		15541 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		15546 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		15557 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		15566 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		15568 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		15570 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		15571 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		15579 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		15588 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		15589 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		15596 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		15606 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		15617 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		15646 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		15650 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		15654 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		15657 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		15664 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		15666 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		15678 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		15679 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		15713 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		15715 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		15723 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		15724 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		15731 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		15737 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		15742 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		15748 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		15759 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		15760 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		15768 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		15772 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		15782 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		15784 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		15830 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		15832 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		15836 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		15845 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		15850 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		15856 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		15861 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		15884 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		15903 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		15909 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		15925 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		15928 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		15929 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		15937 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		15938 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		15947 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		15949 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		15957 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		15964 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		15982 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		15984 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		15996 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		16008 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		16017 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		16020 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		16037 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		16059 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		16081 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		16083 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		16085 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		16102 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		16105 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		16113 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		16114 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		16119 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		16121 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		16132 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		16136 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		16144 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		16146 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		16152 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		16158 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		16165 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		16170 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		16175 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		16176 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		16184 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		16187 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		16190 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		16199 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		16200 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		16216 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		16219 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		16237 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		16242 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		16247 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		16249 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		16254 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		16273 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		16274 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		16282 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		16286 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		16287 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		16302 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		16304 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		16326 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		16327 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		16351 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		16360 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		16363 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		16369 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		16375 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		16380 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		16388 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		16409 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		16412 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		16413 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		16421 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		16442 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		16445 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		16449 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		16459 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		16461 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		16465 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		16468 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		16470 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		16477 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		16483 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		16485 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		16490 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		16491 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		16494 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		16499 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		16506 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		16510 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		16517 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		16534 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		16535 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		16544 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		16557 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		16568 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		16574 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		16585 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		16598 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		16600 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		16603 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		16618 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		16627 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		16632 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		16646 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		16647 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		16654 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		16656 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		16660 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		16662 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		16667 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		16669 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		16677 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		16704 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		16708 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		16717 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		16725 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		16727 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		16732 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		16741 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		16746 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		16748 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		16751 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		16760 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		16765 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		16773 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		16776 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		16789 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		16804 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		16809 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		16815 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		16820 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		16842 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		16855 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		16857 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		16878 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		16879 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		16883 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		16894 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		16906 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		16907 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		16910 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		16913 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		16915 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		16917 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		16919 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		16921 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		16922 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		16925 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		16927 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		16928 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		16929 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		16931 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		16939 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		16948 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		16967 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		16974 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		16977 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		16979 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		16982 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		16987 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		17000 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		17001 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		17003 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		17006 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		17007 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		17013 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		17015 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		17016 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		17017 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		17033 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		17038 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		17055 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		17059 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		17065 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		17067 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		17071 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		17093 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		17096 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		17099 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		17102 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		17109 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		17124 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		17129 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		17141 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		17166 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		17172 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		17184 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		17188 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		17190 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		17191 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		17196 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		17199 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		17207 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		17215 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		17224 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		17229 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		17230 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		17235 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		17243 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		17248 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		17258 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		17259 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		17265 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		17266 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		17279 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		17286 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		17287 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		17294 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		17298 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		17307 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		17318 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		17332 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		17335 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		17340 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		17342 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		17348 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		17353 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		17357 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		17364 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		17378 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		17407 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		17410 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		17437 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		17449 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		17457 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		17469 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		17476 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		17480 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		17501 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		17502 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		17507 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		17510 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		17517 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		17538 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		17540 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		17561 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		17588 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		17589 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		17597 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		17621 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		17626 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		17645 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		17650 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		17667 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		17672 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		17675 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		17690 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		17694 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		17697 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		17698 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		17714 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		17715 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		17724 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		17735 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		17743 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		17745 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		17746 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		17751 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		17760 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		17764 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		17775 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		17778 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		17793 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		17821 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		17824 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		17830 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		17834 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		17835 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		17846 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		17852 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		17853 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		17855 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		17867 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		17878 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		17885 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		17903 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		17904 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		17905 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		17907 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		17908 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		17912 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		17929 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		17937 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		17940 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		17941 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		17947 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		17972 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		17975 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		17976 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		17981 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		17994 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		17995 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		17997 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		18006 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		18007 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		18017 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		18034 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		18044 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		18059 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		18068 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		18079 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		18080 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		18082 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		18083 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		18088 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		18091 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		18093 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		18115 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		18118 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		18122 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		18126 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		18135 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		18153 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		18155 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		18172 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		18194 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		18199 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		18203 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		18222 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		18228 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		18246 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		18260 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		18263 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		18270 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		18278 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		18287 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		18291 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		18293 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		18296 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		18297 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		18303 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		18304 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		18309 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		18310 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		18323 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		18344 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		18346 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		18353 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		18356 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		18377 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		18380 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		18386 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		18389 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		18390 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		18396 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		18398 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		18409 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		18413 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		18416 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		18418 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		18421 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		18423 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		18432 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		18435 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		18436 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		18449 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		18453 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		18460 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		18469 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		18481 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		18489 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		18504 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		18507 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		18511 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		18516 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		18519 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		18524 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		18529 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		18546 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		18550 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		18552 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		18572 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		18574 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		18576 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		18602 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		18603 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		18606 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		18613 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		18626 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		18632 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		18637 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		18638 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		18649 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		18661 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		18666 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		18674 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		18682 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		18707 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		18711 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		18714 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		18719 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		18722 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		18731 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		18738 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		18748 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		18751 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		18753 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		18760 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		18768 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		18770 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		18773 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		18781 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		18782 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		18792 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		18795 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		18826 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		18827 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		18838 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		18844 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		18847 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		18849 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		18858 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		18865 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		18868 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		18870 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		18877 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		18883 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		18887 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		18911 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		18912 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		18939 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		18948 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		18957 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		18958 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		18960 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		18964 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		18965 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		18968 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		18980 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		18984 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		18996 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		18998 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		19027 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		19029 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		19046 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		19048 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		19060 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		19086 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		19122 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		19128 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		19149 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		19154 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		19165 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		19166 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		19170 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		19175 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		19182 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		19183 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		19184 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		19192 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		19204 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		19206 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		19213 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		19217 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		19238 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		19242 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		19243 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		19245 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		19249 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		19252 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		19253 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		19269 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		19281 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		19284 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		19285 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		19287 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		19291 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		19293 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		19296 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		19298 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		19306 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		19313 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		19318 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		19331 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		19336 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		19349 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		19354 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		19355 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		19372 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		19381 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		19382 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		19385 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		19393 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		19406 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		19411 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		19412 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		19414 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		19416 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		19423 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		19430 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		19435 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		19447 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		19453 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		19462 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		19477 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		19487 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		19490 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		19492 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		19494 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		19498 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		19504 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		19508 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		19513 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		19514 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		19517 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		19519 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		19520 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		19528 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		19537 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		19545 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		19557 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		19559 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		19563 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		19564 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		19566 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		19568 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		19570 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		19577 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		19584 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		19585 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		19588 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		19592 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		19609 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		19612 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		19620 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		19669 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		19670 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		19672 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		19676 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		19687 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		19690 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		19691 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		19692 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		19708 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		19711 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		19719 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		19731 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		19734 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		19741 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		19760 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		19762 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		19774 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		19782 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		19784 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		19789 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		19792 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		19811 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		19812 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		19820 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		19822 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		19831 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		19832 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		19836 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		19837 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		19854 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		19867 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		19877 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		19879 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		19885 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		19902 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		19919 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		19921 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		19928 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		19932 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		19935 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		19939 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		19941 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		19952 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		19968 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		19974 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		19985 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		20001 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		20020 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		20027 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		20034 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		20042 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		20051 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		20054 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		20055 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		20061 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		20074 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		20077 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		20080 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		20088 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		20104 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		20105 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		20126 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		20131 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		20157 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		20161 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		20162 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		20165 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		20174 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		20181 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		20182 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		20184 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		20208 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		20210 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		20213 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		20228 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		20248 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		20252 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		20266 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		20292 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		20295 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		20296 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		20297 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		20299 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		20300 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		20311 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		20313 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		20318 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		20324 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		20346 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		20356 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		20372 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		20382 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		20383 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		20386 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		20389 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		20402 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		20418 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		20426 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		20428 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		20431 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		20432 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		20440 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		20447 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		20451 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		20459 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		20460 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		20461 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		20466 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		20468 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		20489 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		20497 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		20504 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		20514 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		20526 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		20527 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		20540 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		20560 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		20561 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		20565 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		20568 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		20573 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		20581 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		20587 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		20594 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		20595 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		20596 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		20597 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		20603 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		20629 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		20630 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		20633 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		20651 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		20669 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		20671 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		20685 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		20694 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		20695 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		20705 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		20706 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		20718 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		20721 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		20722 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		20739 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		20745 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		20754 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		20756 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		20758 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		20763 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		20787 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		20788 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		20801 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		20802 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		20812 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		20815 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		20831 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		20845 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		20856 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		20860 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		20863 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		20865 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		20867 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		20871 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		20876 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		20894 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		20895 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		20905 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		20906 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		20911 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		20953 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		20976 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		20986 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		20989 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		20994 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		21005 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		21008 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		21009 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		21010 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		21020 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		21023 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		21030 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		21035 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		21038 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		21040 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		21042 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		21044 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		21055 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		21068 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		21076 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		21093 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		21102 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		21103 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		21111 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		21119 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		21126 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		21127 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		21130 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		21131 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		21139 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		21142 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		21144 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		21153 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		21157 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		21167 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		21172 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		21176 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		21179 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		21185 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		21195 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		21197 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		21199 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		21202 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		21204 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		21206 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		21211 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		21214 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		21218 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		21225 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		21233 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		21235 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		21237 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		21244 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		21261 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		21272 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		21289 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		21295 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		21296 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		21297 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		21300 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		21303 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		21309 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		21315 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		21318 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		21323 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		21326 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		21327 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		21337 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		21350 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		21352 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		21353 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		21355 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		21359 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		21366 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		21376 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		21377 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		21384 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		21390 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		21397 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		21401 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		21406 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		21409 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		21410 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		21417 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		21419 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		21422 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		21427 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		21431 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		21434 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		21442 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		21443 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		21444 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		21457 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		21468 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		21475 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		21485 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		21495 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		21505 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		21510 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		21513 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		21514 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		21522 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		21524 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		21527 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		21536 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		21541 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		21556 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		21561 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		21576 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		21580 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		21588 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		21598 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		21599 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		21612 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		21619 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		21625 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		21628 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		21661 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		21664 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		21672 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		21677 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		21702 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		21707 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		21709 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		21711 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		21723 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		21729 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		21736 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		21797 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		21802 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		21819 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		21825 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		21829 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		21835 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		21847 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		21849 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		21851 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		21859 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		21862 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		21883 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		21884 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		21886 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		21902 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		21904 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		21905 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		21907 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		21932 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		21935 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		21937 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		21982 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		21997 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		21998 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		22004 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		22005 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		22007 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		22016 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		22017 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		22026 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		22036 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		22043 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		22076 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		22086 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		22094 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		22105 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		22106 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		22107 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		22117 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		22121 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		22123 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		22129 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		22137 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		22141 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		22144 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		22163 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		22169 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		22173 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		22187 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		22189 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		22201 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		22204 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		22207 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		22218 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		22228 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		22233 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		22238 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		22255 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		22267 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		22317 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		22318 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		22321 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		22324 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		22341 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		22344 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		22347 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		22353 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		22356 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		22358 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		22363 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		22367 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		22376 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		22377 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		22390 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		22397 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		22400 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		22432 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		22439 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		22444 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		22460 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		22462 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		22466 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		22470 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		22472 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		22473 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		22474 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		22496 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		22507 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		22509 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		22516 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		22518 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		22529 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		22531 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		22533 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		22535 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		22536 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		22551 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		22554 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		22555 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		22557 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		22562 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		22594 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		22596 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		22609 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		22627 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		22630 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		22634 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		22644 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		22647 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		22652 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		22653 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		22662 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		22668 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		22677 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		22680 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		22711 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		22724 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		22735 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		22738 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		22757 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		22758 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		22770 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		22776 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		22779 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		22780 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		22787 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		22788 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		22789 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		22796 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		22800 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		22803 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		22807 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		22816 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		22820 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		22835 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		22836 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		22844 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		22852 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		22857 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		22865 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		22868 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		22869 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		22872 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		22874 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		22883 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		22896 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		22898 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		22904 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		22913 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		22915 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		22919 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		22922 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		22924 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		22925 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		22927 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		22941 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		22949 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		22950 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		22954 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		22957 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		22972 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		22974 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		22995 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		22996 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		22999 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		23000 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		23005 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		23006 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		23008 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		23017 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		23020 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		23032 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		23042 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		23043 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		23045 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		23053 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		23055 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		23056 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		23059 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		23065 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		23068 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		23073 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		23082 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		23083 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		23089 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		23090 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		23093 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		23096 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		23097 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		23110 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		23112 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		23117 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		23119 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		23121 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		23127 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		23131 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		23137 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		23147 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		23163 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		23166 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		23170 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		23175 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		23190 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		23196 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		23199 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		23201 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		23207 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		23211 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		23214 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		23223 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		23235 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		23237 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		23238 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		23240 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		23243 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		23254 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		23265 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		23274 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		23283 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		23294 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		23296 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		23304 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		23311 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		23327 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		23339 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		23345 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		23355 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		23357 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		23359 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		23365 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		23367 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		23372 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		23382 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		23383 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		23394 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		23397 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		23407 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		23417 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		23419 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		23430 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		23433 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		23436 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		23439 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		23447 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		23453 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		23465 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		23466 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		23472 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		23476 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		23480 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		23483 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		23484 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		23488 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		23491 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		23499 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		23500 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		23502 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		23511 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		23520 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		23529 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		23532 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		23545 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		23548 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		23555 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		23559 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		23560 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		23562 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		23575 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		23585 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		23593 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		23599 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		23610 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		23622 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		23627 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		23654 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		23655 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		23663 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		23668 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		23677 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		23681 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		23695 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		23696 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		23720 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		23733 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		23769 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		23775 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		23793 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		23795 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		23800 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		23822 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		23832 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		23835 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		23840 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		23859 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		23866 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		23873 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		23886 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		23889 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		23891 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		23911 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		23915 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		23917 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		23920 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		23937 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		23941 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		23954 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		23972 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		23975 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		23978 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		23988 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		23992 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		24003 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		24012 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		24016 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		24025 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		24030 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		24034 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		24042 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		24053 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		24066 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		24069 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		24079 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		24081 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		24093 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		24115 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		24133 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		24136 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		24141 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		24157 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		24158 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		24167 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		24178 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		24179 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		24186 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		24188 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		24193 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		24197 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		24201 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		24214 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		24219 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		24244 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		24253 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		24259 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		24261 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		24283 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		24284 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		24294 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		24295 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		24297 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		24298 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		24304 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		24309 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		24328 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		24332 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		24334 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		24339 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		24357 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		24374 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		24387 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		24403 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		24405 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		24417 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		24421 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		24448 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		24465 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		24468 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		24469 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		24473 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		24474 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		24493 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		24496 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		24515 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		24517 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		24522 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		24541 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		24544 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		24548 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		24549 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		24551 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		24553 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		24567 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		24577 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		24593 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		24596 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		24612 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		24613 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		24616 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		24617 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		24630 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		24631 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		24636 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		24637 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		24643 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		24645 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		24646 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		24659 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		24663 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		24686 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		24688 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		24690 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		24705 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		24708 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		24714 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		24715 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		24716 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		24723 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		24735 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		24741 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		24742 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		24746 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		24757 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		24759 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		24770 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		24776 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		24800 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		24818 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		24828 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		24834 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		24837 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		24843 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		24849 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		24863 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		24876 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		24877 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		24878 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		24879 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		24881 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		24893 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		24899 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		24901 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		24902 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		24911 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		24916 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		24918 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		24921 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		24928 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		24937 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		24960 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		24962 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		24964 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		24966 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		24967 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		24995 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		25000 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		25009 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		25013 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		25026 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		25044 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		25083 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		25085 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		25096 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		25099 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		25103 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		25134 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		25139 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		25154 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		25164 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		25173 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		25175 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		25181 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		25183 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		25191 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		25200 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		25210 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		25218 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		25232 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		25247 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		25250 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		25254 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		25258 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		25260 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		25262 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		25265 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		25274 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		25289 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		25292 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		25300 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		25304 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		25308 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		25324 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		25332 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		25333 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		25335 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		25336 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		25344 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		25348 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		25350 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		25354 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		25357 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		25377 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		25378 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		25385 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		25393 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		25395 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		25402 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		25409 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		25411 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		25421 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		25426 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		25433 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		25441 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		25446 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		25457 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		25464 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		25475 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		25479 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		25495 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		25498 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		25504 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		25510 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		25513 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		25525 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		25533 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		25535 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		25549 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		25555 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		25561 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		25568 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		25588 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		25590 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		25604 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		25613 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		25615 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		25617 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		25620 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		25622 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		25624 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		25633 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		25634 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		25645 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		25647 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		25653 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		25658 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		25667 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		25669 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		25671 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		25674 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		25678 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		25684 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		25687 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		25689 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		25695 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		25718 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		25742 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		25744 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		25746 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		25765 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		25771 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		25772 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		25785 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		25790 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		25795 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		25797 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		25798 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		25808 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		25830 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		25854 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		25858 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		25859 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		25865 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		25873 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		25874 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		25881 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		25886 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		25892 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		25906 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		25910 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		25911 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		25941 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		25948 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		25949 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		25972 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		25976 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		25982 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		25995 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		26007 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		26011 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		26027 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		26028 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		26032 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		26038 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		26045 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		26053 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		26054 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		26058 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		26059 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		26061 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		26066 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		26070 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		26073 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		26077 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		26089 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		26093 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		26100 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		26120 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		26139 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		26146 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		26151 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		26158 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		26166 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		26170 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		26172 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		26183 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		26190 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		26195 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		26215 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		26218 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		26220 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		26225 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		26227 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		26231 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		26240 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		26247 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		26248 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		26258 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		26265 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		26266 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		26281 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		26282 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		26292 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		26293 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		26294 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		26299 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		26301 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		26315 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		26325 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		26328 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		26344 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		26346 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		26369 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		26379 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		26387 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		26397 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		26400 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		26402 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		26403 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		26405 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		26413 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		26431 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		26435 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		26438 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		26441 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		26445 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		26454 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		26455 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		26458 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		26466 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		26474 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		26475 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		26477 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		26489 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		26490 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		26492 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		26503 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		26517 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		26519 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		26531 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		26540 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		26545 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		26550 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		26553 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		26560 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		26562 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		26575 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		26576 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		26578 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		26581 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		26589 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		26591 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		26597 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		26599 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		26608 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		26614 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		26617 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		26624 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		26625 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		26634 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		26637 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		26650 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		26654 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		26658 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		26673 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		26674 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		26678 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		26688 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		26690 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		26691 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		26714 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		26718 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		26721 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		26728 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		26732 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		26734 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		26765 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		26782 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		26784 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		26797 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		26801 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		26802 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		26804 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		26806 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		26807 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		26812 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		26825 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		26830 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		26835 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		26839 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		26846 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		26862 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		26866 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		26867 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		26870 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		26876 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		26883 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		26903 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		26906 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		26926 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		26931 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		26940 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		26959 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		26964 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		26970 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		26982 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		26986 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		27003 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		27010 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		27011 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		27041 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		27044 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		27053 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		27055 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		27086 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		27096 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		27101 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		27104 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		27116 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		27128 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		27133 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		27134 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		27140 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		27151 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		27160 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		27175 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		27177 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		27188 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		27197 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		27208 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		27209 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		27227 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		27245 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		27247 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		27259 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		27286 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		27294 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		27317 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		27318 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		27338 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		27342 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		27359 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		27366 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		27376 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		27377 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		27382 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		27388 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		27398 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		27400 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		27406 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		27407 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		27414 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		27416 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		27419 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		27422 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		27442 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		27452 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		27461 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		27463 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		27490 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		27492 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		27497 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		27510 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		27513 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		27514 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		27524 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		27540 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		27542 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		27560 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		27569 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		27572 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		27573 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		27575 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		27584 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		27597 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		27599 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		27605 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		27613 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		27623 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		27630 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		27637 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		27644 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		27650 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		27664 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		27670 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		27677 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		27678 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		27695 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		27696 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		27701 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		27707 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		27708 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		27711 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		27713 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		27715 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		27719 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		27723 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		27726 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		27738 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		27752 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		27761 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		27763 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		27766 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		27777 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		27778 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		27786 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		27788 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		27804 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		27808 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		27813 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		27834 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		27852 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		27853 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		27872 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		27874 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		27893 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		27901 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		27902 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		27909 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		27910 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		27914 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		27920 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		27922 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		27933 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		27939 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		27942 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		27946 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		27948 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		27949 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		27953 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		27954 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		27961 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		27965 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		27969 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		27971 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		27977 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		27978 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		27984 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		27991 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		27994 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		27995 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		28002 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		28004 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		28005 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		28006 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		28010 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		28020 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		28021 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		28033 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		28036 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		28047 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		28054 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		28064 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		28073 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		28080 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		28090 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		28093 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		28097 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		28114 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		28115 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		28132 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		28142 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		28143 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		28164 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		28167 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		28169 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		28172 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		28175 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		28185 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		28193 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		28196 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		28211 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		28225 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		28228 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		28233 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		28242 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		28244 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		28255 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		28259 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		28261 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		28284 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		28287 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		28290 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		28293 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		28302 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		28308 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		28321 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		28323 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		28330 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		28340 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		28359 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		28379 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		28381 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		28382 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		28397 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		28406 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		28415 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		28417 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		28422 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		28447 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		28460 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		28466 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		28467 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		28491 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		28500 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		28507 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		28512 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		28515 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		28517 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		28521 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		28525 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		28527 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		28529 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		28530 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		28533 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		28539 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		28540 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		28558 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		28563 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		28580 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		28589 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		28602 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		28608 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		28619 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		28620 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		28644 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		28646 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		28650 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		28652 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		28666 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		28669 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		28673 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		28679 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		28683 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		28690 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		28698 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		28702 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		28714 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		28728 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		28733 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		28738 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		28743 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		28767 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		28773 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		28775 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		28776 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		28783 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		28797 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		28805 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		28806 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		28812 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		28816 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		28831 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		28847 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		28859 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		28860 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		28868 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		28871 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		28874 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		28878 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		28885 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		28897 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		28902 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		28913 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		28915 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		28934 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		28961 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		28968 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		28978 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		28986 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		28993 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		28995 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		28998 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		29005 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		29019 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		29020 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		29024 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		29041 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		29048 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		29052 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		29053 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		29055 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		29060 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		29073 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		29075 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		29082 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		29084 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		29086 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		29087 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		29096 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		29100 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		29105 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		29122 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		29140 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		29141 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		29150 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		29154 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		29164 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		29168 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		29170 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		29175 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		29184 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		29187 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		29198 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		29204 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		29207 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		29211 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		29219 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		29223 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		29227 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		29229 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		29234 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		29235 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		29238 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		29241 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		29243 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		29249 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		29254 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		29256 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		29285 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		29305 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		29313 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		29316 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		29325 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		29327 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		29334 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		29335 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		29342 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		29348 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		29354 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		29363 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		29365 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		29369 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		29371 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		29372 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		29375 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		29379 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		29386 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		29403 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		29407 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		29408 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		29409 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		29413 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		29424 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		29430 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		29432 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		29436 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		29442 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		29446 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		29448 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		29451 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		29470 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		29471 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		29475 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		29492 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		29503 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		29504 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		29512 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		29517 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		29527 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		29529 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		29531 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		29539 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		29541 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		29552 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		29560 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		29569 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		29570 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		29581 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		29588 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		29604 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		29610 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		29625 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		29641 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		29649 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		29655 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		29656 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		29660 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		29690 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		29704 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		29709 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		29712 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		29716 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		29725 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		29735 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		29737 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		29782 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		29791 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		29793 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		29804 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		29816 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		29826 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		29828 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		29846 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		29849 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		29853 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		29872 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		29885 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		29891 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		29904 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		29911 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		29914 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		29915 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		29922 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		29924 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		29926 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		29929 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		29943 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		29946 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		29947 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		29949 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		29950 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		29983 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		29989 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		29990 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		29991 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		29996 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		29999 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		30014 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		30016 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		30020 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		30028 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		30029 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		30036 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		30041 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		30045 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		30046 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		30047 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		30053 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		30055 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		30064 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		30068 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		30074 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		30081 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		30084 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		30090 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		30107 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		30109 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		30112 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		30117 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		30139 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		30154 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		30171 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		30189 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		30190 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		30191 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		30192 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		30208 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		30217 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		30234 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		30250 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		30265 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		30267 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		30275 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		30280 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		30290 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		30296 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		30298 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		30302 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		30319 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		30326 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		30344 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		30360 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		30363 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		30374 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		30379 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		30384 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		30385 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		30393 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		30400 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		30409 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		30411 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		30419 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		30420 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		30425 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		30428 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		30429 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		30430 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		30442 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		30445 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		30451 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		30453 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		30457 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		30458 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		30466 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		30470 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		30475 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		30476 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		30477 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		30484 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		30489 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		30500 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		30513 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		30523 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		30536 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		30537 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		30541 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		30545 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		30576 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		30578 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		30580 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		30582 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		30584 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		30585 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		30586 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		30587 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		30591 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		30601 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		30603 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		30612 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		30639 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		30641 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		30644 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		30657 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		30661 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		30679 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		30684 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		30686 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		30695 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		30697 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		30710 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		30712 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		30720 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		30722 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		30725 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		30726 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		30737 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		30738 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		30744 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		30771 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		30781 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		30783 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		30805 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		30807 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		30811 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		30817 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		30829 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		30831 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		30844 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		30860 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		30869 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		30873 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		30890 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		30897 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		30913 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		30923 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		30930 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		30951 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		30965 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		30967 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		30983 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		30987 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		30989 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		30995 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		30997 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		31001 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		31007 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		31010 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		31011 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		31012 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		31031 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		31034 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		31035 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		31038 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		31054 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		31077 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		31080 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		31096 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		31115 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		31135 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		31137 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		31144 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		31157 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		31179 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		31181 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		31190 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		31192 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		31217 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		31218 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		31224 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		31235 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		31248 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		31257 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		31261 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		31272 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		31274 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		31284 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		31291 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		31292 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		31299 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		31303 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		31309 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		31313 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		31315 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		31316 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		31322 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		31331 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		31333 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		31334 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		31336 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		31341 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		31344 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		31348 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		31356 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		31363 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		31383 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		31393 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		31399 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		31403 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		31404 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		31417 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		31418 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		31421 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		31442 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		31457 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		31466 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		31468 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		31474 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		31480 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		31488 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		31490 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		31497 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		31519 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		31525 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		31534 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		31544 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		31560 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		31574 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		31579 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		31591 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		31593 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		31604 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		31617 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		31618 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		31636 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		31645 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		31649 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		31654 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		31666 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		31675 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		31680 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		31686 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		31693 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		31706 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		31713 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		31714 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		31718 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		31721 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		31724 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		31737 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		31741 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		31747 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		31759 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		31764 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		31775 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		31795 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		31835 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		31837 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		31841 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		31842 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		31850 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		31852 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		31857 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		31862 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		31879 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		31889 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		31891 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		31901 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		31912 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		31913 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		31919 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		31922 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		31934 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		31937 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		31941 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		31952 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		31963 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		31968 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		31969 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		31971 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		31974 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		31978 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		31987 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		31999 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		32004 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		32011 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		32016 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		32077 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		32097 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		32110 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		32118 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		32130 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		32131 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		32143 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		32145 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		32152 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		32176 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		32177 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		32182 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		32183 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		32188 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		32201 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		32217 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		32225 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		32234 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		32238 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		32247 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		32254 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		32255 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		32258 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		32262 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		32265 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		32268 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		32269 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		32296 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		32298 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		32299 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		32307 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		32308 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		32314 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		32324 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		32332 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		32333 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		32343 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		32347 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		32352 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		32358 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		32359 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		32364 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		32367 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		32368 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		32370 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		32376 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		32377 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		32385 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		32386 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		32389 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		32398 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		32404 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		32406 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		32407 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		32409 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		32418 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		32420 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		32425 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		32428 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		32430 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		32433 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		32438 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		32462 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		32469 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		32477 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		32501 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		32506 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		32514 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		32528 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		32533 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		32540 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		32541 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		32545 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		32549 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		32552 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		32555 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		32561 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		32571 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		32579 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		32587 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		32588 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		32589 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		32602 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		32614 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		32621 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		32630 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		32640 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		32641 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		32651 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		32652 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		32670 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		32687 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		32711 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		32715 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		32719 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		32722 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		32729 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		32735 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		32736 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		32741 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		32742 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		32745 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		32759 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		32765 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		32768 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		32770 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		32776 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		32777 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		32793 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		32795 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		32796 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		32800 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		32803 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		32807 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		32814 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		32815 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		32820 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		32833 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		32835 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		32846 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		32850 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		32855 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		32856 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		32860 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		32869 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		32876 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		32885 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		32888 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		32890 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		32896 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		32902 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		32904 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		32918 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		32925 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		32939 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		32941 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		32958 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		32989 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		32994 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		33002 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		33007 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		33016 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		33039 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		33041 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		33059 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		33066 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		33071 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		33086 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		33087 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		33088 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		33093 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		33094 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		33107 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		33108 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		33131 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		33132 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		33133 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		33149 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		33151 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		33158 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		33164 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		33165 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		33181 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		33186 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		33190 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		33191 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		33193 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		33194 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		33200 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		33229 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		33232 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		33235 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		33238 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		33242 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		33245 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		33246 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		33248 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		33254 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		33256 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		33270 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		33276 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		33283 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		33297 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		33301 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		33304 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		33309 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		33311 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		33312 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		33313 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		33314 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		33315 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		33318 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		33320 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		33350 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		33369 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		33370 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		33374 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		33376 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		33387 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		33390 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		33403 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		33409 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		33428 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		33432 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		33438 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		33450 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		33457 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		33463 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		33466 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		33470 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		33474 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		33478 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		33484 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		33490 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		33496 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		33502 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		33509 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		33519 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		33536 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		33540 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		33542 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		33546 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		33569 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		33581 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		33588 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		33589 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		33590 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		33595 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		33601 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		33611 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		33621 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		33622 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		33630 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		33642 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		33645 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		33646 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		33649 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		33654 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		33655 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		33663 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		33669 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		33676 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		33679 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		33686 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		33689 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		33703 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		33706 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		33714 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		33716 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		33719 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		33734 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		33743 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		33750 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		33766 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		33769 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		33776 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		33785 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		33786 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		33787 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		33812 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		33822 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		33826 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		33831 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		33841 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		33849 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		33856 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		33857 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		33864 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		33866 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		33879 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		33885 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		33889 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		33893 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		33905 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		33906 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		33908 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		33909 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		33915 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		33917 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		33936 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		33940 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		33941 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		33950 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		33952 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		33954 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		33957 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		33961 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		33972 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		33973 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		33985 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		33988 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		33996 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		34001 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		34003 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		34013 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		34019 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		34024 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		34038 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		34041 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		34043 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		34051 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		34055 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		34062 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		34067 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		34075 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		34076 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		34078 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		34090 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		34095 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		34098 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		34109 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		34116 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		34122 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		34123 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		34127 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		34128 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		34129 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		34130 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		34133 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		34136 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		34140 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		34147 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		34163 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		34165 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		34171 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		34176 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		34180 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		34183 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		34191 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		34197 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		34213 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		34219 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		34220 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		34223 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		34225 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		34230 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		34231 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		34232 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		34243 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		34277 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		34283 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		34292 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		34293 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		34306 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		34320 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		34330 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		34334 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		34353 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		34359 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		34362 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		34370 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		34380 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		34385 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		34386 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		34390 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		34395 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		34396 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		34400 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		34402 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		34406 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		34407 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		34408 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		34409 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		34411 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		34413 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		34420 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		34425 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		34426 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		34434 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		34435 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		34436 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		34440 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		34448 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		34459 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		34464 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		34469 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		34488 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		34490 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		34496 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		34497 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		34501 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		34507 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		34517 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		34519 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		34523 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		34535 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		34538 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		34544 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		34547 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		34548 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		34559 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		34560 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		34568 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		34579 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		34583 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		34585 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		34615 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		34630 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		34634 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		34645 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		34652 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		34654 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		34655 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		34664 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		34671 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		34673 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		34675 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		34676 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		34678 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		34679 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		34688 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		34689 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		34696 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		34703 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		34730 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		34745 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		34747 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		34751 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		34757 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		34830 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		34833 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		34845 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		34851 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		34858 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		34861 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		34865 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		34871 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		34874 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		34875 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		34884 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		34890 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		34892 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		34910 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		34918 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		34926 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		34927 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		34930 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		34932 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		34952 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		34953 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		34965 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		34970 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		34983 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		34987 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		34991 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		34993 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		35008 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		35010 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		35017 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		35020 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		35022 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		35031 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		35050 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		35051 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		35053 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		35057 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		35059 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		35064 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		35080 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		35087 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		35095 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		35105 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		35113 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		35114 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		35116 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		35134 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		35137 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		35144 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		35160 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		35163 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		35172 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		35179 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		35186 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		35194 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		35207 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		35221 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		35225 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		35227 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		35228 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		35239 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		35246 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		35248 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		35250 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		35264 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		35265 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		35270 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		35277 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		35285 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		35291 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		35297 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		35298 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		35300 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		35301 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		35307 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		35312 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		35316 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		35321 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		35327 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		35331 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		35349 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		35353 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		35365 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		35370 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		35375 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		35387 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		35406 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		35428 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		35431 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		35435 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		35437 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		35438 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		35442 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		35454 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		35462 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		35464 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		35473 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		35484 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		35490 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		35496 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		35505 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		35527 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		35534 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		35535 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		35536 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		35538 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		35545 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		35551 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		35571 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		35578 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		35595 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		35597 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		35599 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		35629 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		35640 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		35645 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		35646 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		35653 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		35655 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		35660 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		35661 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		35669 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		35671 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		35680 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		35681 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		35685 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		35686 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		35687 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		35693 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		35698 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		35700 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		35703 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		35705 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		35710 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		35714 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		35721 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		35723 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		35736 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		35746 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		35770 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		35779 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		35786 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		35792 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		35794 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		35802 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		35810 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		35813 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		35821 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		35827 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		35831 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		35836 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		35838 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		35842 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		35844 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		35847 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		35887 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		35898 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		35916 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		35922 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		35926 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		35942 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		35955 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		35958 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		35965 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		35971 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		35972 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		35979 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		35986 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		35989 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		35995 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		36002 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		36009 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		36016 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		36032 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		36033 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		36037 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		36046 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		36058 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		36064 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		36072 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		36077 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		36079 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		36082 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		36086 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		36089 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		36096 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		36101 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		36111 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		36115 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		36127 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		36128 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		36134 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		36138 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		36140 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		36144 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		36151 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		36155 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		36157 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		36159 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		36161 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		36170 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		36180 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		36186 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		36189 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		36191 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		36207 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		36223 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		36230 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		36231 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		36292 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		36302 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		36303 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		36309 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		36315 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		36322 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		36326 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		36329 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		36333 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		36335 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		36336 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		36338 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		36339 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		36346 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		36364 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		36365 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		36369 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		36370 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		36391 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		36398 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		36402 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		36407 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		36412 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		36422 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		36432 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		36433 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		36443 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		36454 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		36458 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		36459 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		36464 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		36479 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		36501 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		36511 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		36514 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		36516 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		36522 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		36530 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		36539 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		36562 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		36566 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		36568 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		36571 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		36580 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		36585 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		36589 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		36592 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		36593 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		36597 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		36599 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		36600 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		36602 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		36605 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		36607 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		36612 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		36617 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		36619 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		36622 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		36630 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		36635 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		36642 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		36651 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		36663 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		36667 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		36671 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		36693 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		36706 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		36707 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		36714 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		36718 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		36725 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		36727 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		36731 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		36734 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		36741 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		36745 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		36753 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		36766 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		36770 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		36777 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		36786 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		36789 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		36790 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		36791 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		36795 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		36796 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		36807 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		36809 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		36818 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		36819 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		36827 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		36831 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		36832 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		36854 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		36866 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		36895 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		36896 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		36897 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		36900 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		36917 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		36918 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		36920 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		36926 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		36929 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		36933 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		36946 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		36954 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		36955 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		36957 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		36958 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		36967 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		36969 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		36977 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		36978 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		36988 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		36992 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		36994 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		36995 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		37002 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		37004 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		37006 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		37007 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		37015 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		37016 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		37017 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		37019 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		37024 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		37025 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		37026 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		37037 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		37041 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		37053 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		37058 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		37062 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		37085 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		37089 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		37098 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		37108 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		37119 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		37126 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		37134 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		37151 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		37162 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		37168 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		37186 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		37189 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		37190 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		37191 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		37192 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		37194 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		37203 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		37205 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		37219 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		37220 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		37221 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		37224 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		37234 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		37246 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		37263 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		37264 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		37269 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		37290 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		37291 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		37298 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		37302 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		37321 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		37332 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		37334 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		37339 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		37355 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		37359 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		37362 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		37368 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		37378 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		37404 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		37416 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		37419 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		37431 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		37434 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		37435 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		37440 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		37447 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		37463 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		37464 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		37487 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		37490 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		37493 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		37494 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		37504 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		37505 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		37519 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		37520 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		37522 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		37523 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		37531 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		37536 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		37537 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		37542 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		37545 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		37547 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		37563 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		37567 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		37569 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		37572 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		37578 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		37583 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		37598 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		37601 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		37607 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		37609 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		37616 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		37623 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		37626 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		37629 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		37637 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		37643 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		37645 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		37651 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		37654 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		37655 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		37660 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		37669 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		37674 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		37676 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		37690 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		37697 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		37704 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		37706 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		37711 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		37720 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		37734 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		37737 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		37754 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		37766 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		37767 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		37790 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		37803 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		37812 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		37816 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		37836 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		37852 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		37859 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		37864 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		37871 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		37872 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		37873 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		37887 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		37890 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		37892 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		37897 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		37901 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		37903 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		37905 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		37918 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		37923 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		37927 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		37941 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		37949 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		37951 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		37971 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		37973 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		37976 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		37977 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		37981 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		38009 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		38016 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		38029 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		38034 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		38039 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		38042 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		38044 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		38058 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		38061 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		38065 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		38068 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		38079 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		38088 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		38090 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		38097 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		38101 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		38118 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		38126 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		38154 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		38162 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		38164 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		38187 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		38189 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		38190 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		38191 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		38210 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		38217 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		38221 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		38222 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		38225 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		38228 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		38229 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		38241 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		38242 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		38243 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		38249 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		38251 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		38259 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		38264 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		38267 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		38274 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		38278 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		38289 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		38320 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		38334 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		38350 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		38352 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		38364 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		38392 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		38403 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		38406 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		38415 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		38431 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		38446 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		38454 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		38465 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		38471 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		38477 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		38484 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		38490 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		38492 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		38505 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		38511 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		38514 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		38517 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		38533 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		38543 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		38551 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		38552 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		38557 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		38568 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		38573 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		38576 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		38589 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		38604 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		38606 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		38612 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		38615 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		38616 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		38619 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		38622 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		38633 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		38646 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		38655 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		38656 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		38661 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		38663 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		38666 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		38672 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		38683 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		38692 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		38699 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		38700 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		38701 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		38706 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		38718 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		38722 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		38728 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		38731 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		38737 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		38739 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		38742 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		38747 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		38757 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		38760 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		38762 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		38772 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		38782 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		38785 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		38787 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		38801 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		38814 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		38821 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		38837 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		38848 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		38858 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		38860 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		38872 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		38882 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		38884 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		38897 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		38901 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		38903 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		38905 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		38907 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		38908 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		38924 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		38935 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		38938 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		38941 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		38945 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		38948 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		38952 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		38956 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		38957 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		38958 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		38960 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		38961 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		38965 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		38968 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		38971 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		38972 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		38975 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		38996 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		39003 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		39010 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		39034 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		39046 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		39051 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		39052 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		39053 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		39054 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		39055 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		39057 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		39064 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		39065 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		39076 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		39101 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		39111 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		39115 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		39121 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		39122 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		39124 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		39125 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		39128 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		39133 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		39139 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		39153 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		39154 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		39155 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		39161 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		39163 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		39171 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		39174 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		39180 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		39181 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		39184 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		39197 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		39221 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		39227 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		39248 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		39252 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		39264 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		39280 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		39282 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		39285 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		39287 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		39295 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		39303 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		39316 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		39318 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		39332 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		39333 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		39346 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		39348 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		39351 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		39355 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		39361 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		39371 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		39388 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		39414 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		39416 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		39421 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		39430 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		39433 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		39448 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		39450 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		39455 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		39456 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		39461 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		39474 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		39475 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		39482 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		39487 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		39488 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		39496 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		39506 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		39520 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		39522 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		39536 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		39544 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		39550 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		39558 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		39562 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		39584 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		39590 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		39594 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		39600 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		39606 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		39609 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		39614 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		39624 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		39630 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		39634 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		39635 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		39639 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		39643 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		39646 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		39655 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		39656 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		39672 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		39680 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		39681 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		39682 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		39691 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		39707 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		39711 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		39712 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		39716 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		39727 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		39732 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		39734 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		39744 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		39750 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		39754 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		39771 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		39783 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		39793 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		39805 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		39811 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		39813 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		39816 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		39819 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		39839 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		39842 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		39855 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		39858 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		39859 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		39879 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		39896 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		39902 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		39914 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		39917 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		39930 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		39936 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		39945 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		39959 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		39962 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		39968 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		39971 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		39975 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		39995 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		40004 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		40008 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		40009 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		40010 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		40013 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		40016 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		40036 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		40038 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		40059 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		40064 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		40068 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		40074 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		40084 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		40098 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		40106 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		40110 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		40113 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		40126 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		40131 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		40140 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		40141 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		40158 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		40165 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		40171 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		40177 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		40178 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		40187 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		40196 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		40202 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		40229 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		40231 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		40241 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		40251 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		40255 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		40256 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		40277 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		40278 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		40288 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		40291 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		40294 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		40303 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		40324 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		40327 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		40333 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		40346 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		40369 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		40370 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		40377 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		40378 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		40382 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		40392 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		40404 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		40407 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		40422 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		40429 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		40431 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		40436 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		40445 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		40447 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		40464 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		40471 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		40473 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		40475 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		40485 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		40486 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		40498 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		40500 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		40509 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		40511 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		40532 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		40542 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		40545 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		40547 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		40555 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		40577 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		40579 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		40601 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		40628 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		40629 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		40630 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		40635 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		40636 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		40638 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		40641 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		40653 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		40658 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		40659 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		40660 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		40661 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		40667 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		40678 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		40685 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		40694 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		40696 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		40698 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		40699 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		40704 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		40720 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		40724 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		40757 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		40767 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		40772 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		40780 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		40785 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		40792 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		40793 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		40794 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		40810 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		40819 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		40827 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		40833 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		40873 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		40877 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		40878 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		40887 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		40891 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		40901 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		40902 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		40905 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		40907 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		40909 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		40910 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		40931 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		40943 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		40964 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		40966 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		40968 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		40969 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		40972 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		40976 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		40984 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		40999 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		41002 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		41006 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		41029 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		41055 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		41060 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		41066 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		41068 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		41070 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		41079 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		41082 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		41084 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		41113 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		41115 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		41120 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		41122 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		41138 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		41141 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		41144 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		41146 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		41153 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		41156 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		41157 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		41165 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		41169 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		41191 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		41193 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		41195 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		41196 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		41215 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		41219 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		41222 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		41233 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		41252 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		41262 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		41276 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		41285 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		41294 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		41301 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		41308 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		41319 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		41327 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		41328 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		41330 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		41336 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		41339 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		41344 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		41376 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		41387 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		41391 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		41397 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		41401 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		41408 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		41413 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		41434 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		41437 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		41440 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		41460 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		41464 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		41470 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		41480 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		41509 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		41514 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		41526 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		41531 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		41545 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		41554 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		41562 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		41566 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		41570 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		41579 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		41584 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		41593 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		41627 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		41629 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		41632 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		41647 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		41651 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		41653 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		41659 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		41667 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		41671 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		41673 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		41677 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		41685 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		41690 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		41691 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		41695 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		41710 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		41745 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		41750 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		41752 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		41754 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		41765 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		41767 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		41804 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		41805 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		41807 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		41808 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		41828 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		41830 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		41832 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		41835 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		41845 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		41849 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		41852 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		41853 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		41856 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		41859 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		41861 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		41872 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		41873 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		41877 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		41904 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		41909 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		41912 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		41923 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		41931 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		41946 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		41952 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		41955 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		41962 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		41974 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		41979 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		41981 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		41986 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		41994 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		42000 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		42005 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		42014 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		42019 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		42020 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		42024 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		42027 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		42040 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		42041 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		42045 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		42050 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		42061 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		42069 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		42071 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		42094 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		42105 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		42112 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		42113 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		42132 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		42145 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		42156 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		42169 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		42187 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		42189 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		42207 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		42215 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		42221 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		42237 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		42239 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		42247 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		42249 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		42250 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		42253 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		42262 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		42266 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		42268 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		42290 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		42298 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		42319 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		42347 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		42354 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		42365 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		42370 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		42372 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		42380 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		42387 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		42397 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		42398 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		42400 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		42401 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		42403 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		42405 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		42428 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		42429 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		42430 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		42431 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		42436 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		42439 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		42444 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		42445 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		42448 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		42454 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		42473 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		42483 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		42485 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		42495 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		42513 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		42514 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		42517 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		42525 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		42527 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		42532 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		42534 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		42552 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		42553 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		42555 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		42564 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		42577 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		42582 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		42592 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		42597 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		42599 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		42610 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		42614 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		42619 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		42627 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		42628 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		42630 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		42633 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		42637 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		42673 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		42679 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		42689 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		42702 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		42703 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		42707 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		42714 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		42715 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		42723 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		42729 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		42732 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		42734 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		42739 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		42759 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		42764 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		42769 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		42778 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		42786 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		42792 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		42813 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		42826 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		42827 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		42834 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		42845 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		42849 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		42864 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		42870 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		42878 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		42879 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		42880 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		42881 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		42887 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		42890 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		42898 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		42899 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		42922 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		42927 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		42931 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		42943 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		42946 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		42956 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		42957 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		42962 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		42985 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		42990 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		42991 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		43002 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		43004 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		43005 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		43015 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		43019 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		43029 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		43030 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		43031 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		43041 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		43046 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		43047 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		43048 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		43061 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		43069 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		43074 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		43077 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		43079 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		43084 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		43088 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		43093 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		43098 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		43103 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		43106 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		43118 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		43126 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		43131 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		43132 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		43134 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		43142 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		43152 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		43153 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		43154 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		43164 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		43166 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		43176 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		43179 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		43204 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		43206 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		43208 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		43214 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		43224 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		43229 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		43244 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		43245 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		43248 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		43256 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		43260 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		43263 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		43265 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		43293 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		43300 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		43335 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		43336 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		43341 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		43346 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		43356 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		43361 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		43367 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		43371 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		43385 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		43394 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		43397 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		43403 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		43408 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		43425 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		43437 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		43443 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		43447 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		43450 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		43453 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		43454 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		43461 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		43462 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		43466 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		43479 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		43481 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		43483 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		43485 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		43492 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		43510 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		43511 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		43514 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		43525 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		43527 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		43528 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		43533 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		43544 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		43551 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		43560 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		43566 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		43587 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		43592 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		43595 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		43596 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		43601 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		43613 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		43615 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		43635 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		43638 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		43646 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		43647 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		43661 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		43674 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		43675 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		43680 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		43684 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		43687 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		43688 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		43689 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		43702 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		43709 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		43712 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		43718 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		43723 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		43737 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		43742 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		43757 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		43759 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		43768 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		43771 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		43774 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		43780 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		43781 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		43784 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		43803 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		43810 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		43820 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		43861 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		43863 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		43865 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		43870 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		43876 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		43881 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		43887 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		43888 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		43889 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		43890 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		43895 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		43899 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		43900 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		43916 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		43919 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		43922 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		43927 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		43929 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		43932 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		43933 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		43937 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		43945 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		43947 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		43954 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		43967 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		43979 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		43982 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		43997 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		43999 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		44009 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		44010 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		44017 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		44025 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		44032 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		44038 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		44039 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		44045 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		44053 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		44057 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		44075 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		44076 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		44080 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		44086 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		44088 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		44092 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		44094 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		44097 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		44098 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		44101 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		44106 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		44111 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		44113 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		44128 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		44131 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		44138 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		44141 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		44143 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		44158 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		44171 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		44176 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		44187 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		44189 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		44193 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		44197 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		44209 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		44214 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		44218 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		44219 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		44220 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		44224 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		44229 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		44237 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		44243 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		44244 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		44255 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		44256 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		44262 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		44263 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		44264 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		44268 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		44277 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		44280 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		44283 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		44290 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		44292 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		44297 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		44302 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		44315 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		44334 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		44335 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		44355 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		44364 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		44398 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		44401 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		44406 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		44422 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		44425 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		44426 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		44434 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		44447 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		44477 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		44506 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		44507 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		44510 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		44526 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		44527 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		44535 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		44538 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		44541 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		44549 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		44559 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		44576 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		44580 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		44583 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		44587 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		44598 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		44619 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		44620 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		44650 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		44656 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		44658 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		44659 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		44696 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		44697 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		44709 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		44710 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		44731 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		44737 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		44740 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		44741 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		44742 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		44762 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		44771 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		44788 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		44796 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		44797 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		44805 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		44813 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		44838 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		44840 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		44853 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		44855 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		44856 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		44861 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		44863 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		44866 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		44876 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		44883 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		44884 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		44892 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		44904 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		44910 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		44913 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		44918 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		44926 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		44930 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		44937 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		44943 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		44952 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		44963 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		44974 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		44977 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		44982 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		44988 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		44992 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		45002 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		45006 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		45012 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		45014 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		45019 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		45022 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		45027 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		45039 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		45041 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		45048 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		45064 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		45082 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		45085 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		45095 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		45103 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		45134 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		45144 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		45148 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		45150 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		45153 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		45158 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		45165 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		45177 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		45178 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		45185 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		45201 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		45205 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		45206 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		45221 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		45228 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		45232 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		45239 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		45245 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		45251 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		45254 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		45260 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		45263 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		45265 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		45269 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		45285 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		45302 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		45306 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		45320 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		45330 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		45338 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		45341 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		45343 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		45360 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		45361 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		45364 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		45370 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		45378 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		45389 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		45397 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		45404 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		45409 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		45410 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		45463 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		45472 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		45475 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		45478 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		45491 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		45493 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		45502 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		45503 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		45505 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		45506 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		45514 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		45522 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		45525 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		45531 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		45534 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		45544 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		45550 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		45553 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		45559 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		45574 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		45579 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		45584 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		45591 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		45592 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		45593 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		45599 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		45604 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		45605 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		45609 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		45618 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		45640 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		45641 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		45648 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		45651 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		45652 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		45656 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		45659 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		45663 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		45671 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		45676 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		45677 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		45695 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		45701 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		45705 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		45706 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		45723 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		45735 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		45756 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		45763 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		45771 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		45775 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		45776 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		45778 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		45779 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		45780 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		45786 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		45789 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		45790 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		45793 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		45812 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		45814 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		45829 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		45835 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		45856 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		45857 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		45861 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		45863 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		45879 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		45891 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		45892 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		45897 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		45913 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		45920 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		45927 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		45930 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		45931 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		45938 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		45987 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		45993 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		45995 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		46007 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		46008 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		46012 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		46017 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		46024 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		46026 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		46027 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		46043 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		46049 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		46056 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		46063 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		46065 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		46070 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		46073 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		46078 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		46085 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		46093 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		46104 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		46105 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		46133 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		46136 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		46138 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		46150 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		46162 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		46163 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		46169 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		46175 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		46177 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		46192 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		46195 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		46207 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		46249 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		46253 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		46264 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		46271 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		46278 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		46290 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		46303 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		46308 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		46309 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		46314 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		46318 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		46321 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		46330 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		46342 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		46349 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		46352 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		46379 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		46381 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		46382 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		46386 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		46387 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		46395 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		46407 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		46411 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		46418 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		46420 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		46426 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		46427 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		46431 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		46448 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		46449 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		46466 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		46470 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		46473 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		46492 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		46493 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		46519 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		46524 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		46545 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		46546 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		46550 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		46551 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		46555 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		46559 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		46561 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		46569 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		46575 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		46580 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		46613 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		46614 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		46617 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		46620 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		46622 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		46626 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		46629 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		46638 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		46641 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		46654 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		46662 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		46666 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		46672 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		46678 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		46682 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		46685 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		46689 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		46692 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		46699 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		46704 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		46717 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		46721 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		46726 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		46732 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		46734 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		46744 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		46764 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		46765 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		46768 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		46777 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		46778 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		46781 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		46795 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		46801 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		46810 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		46814 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		46817 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		46818 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		46824 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		46825 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		46831 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		46838 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		46841 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		46868 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		46873 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		46882 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		46903 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		46914 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		46919 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		46921 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		46922 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		46930 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		46937 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		46940 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		46956 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		46958 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		46967 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		46969 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		46970 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		46971 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		46973 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		46980 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		46995 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		47001 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		47014 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		47015 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		47016 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		47018 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		47062 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		47065 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		47070 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		47071 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		47075 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		47076 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		47077 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		47084 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		47087 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		47113 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		47117 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		47122 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		47124 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		47126 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		47131 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		47140 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		47150 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		47160 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		47164 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		47166 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		47167 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		47178 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		47186 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		47187 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		47189 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		47190 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		47194 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		47201 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		47204 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		47218 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		47219 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		47226 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		47230 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		47245 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		47257 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		47260 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		47266 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		47272 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		47290 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		47299 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		47307 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		47317 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		47332 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		47336 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		47355 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		47365 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		47367 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		47379 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		47382 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		47399 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		47401 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		47403 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		47410 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		47421 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		47432 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		47442 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		47451 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		47463 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		47466 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		47467 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		47479 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		47483 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		47484 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		47489 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		47498 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		47499 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		47507 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		47526 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		47534 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		47538 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		47539 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		47544 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		47548 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		47557 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		47564 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		47568 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		47583 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		47584 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		47599 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		47601 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		47614 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		47618 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		47625 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		47626 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		47627 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		47629 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		47635 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		47652 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		47660 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		47665 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		47677 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		47692 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		47703 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		47711 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		47724 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		47734 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		47735 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		47751 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		47768 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		47773 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		47777 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		47780 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		47781 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		47791 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		47793 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		47800 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		47801 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		47807 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		47808 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		47818 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		47834 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		47836 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		47837 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		47848 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		47861 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		47862 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		47864 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		47870 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		47892 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		47906 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		47910 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		47939 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		47944 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		47950 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		47951 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		47952 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		47957 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		47959 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		47964 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		47967 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		47973 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		47987 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		47989 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		48000 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		48021 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		48039 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		48041 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		48046 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		48050 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		48052 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		48053 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		48068 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		48072 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		48073 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		48085 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		48102 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		48104 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		48106 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		48113 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		48122 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		48127 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		48130 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		48131 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		48132 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		48137 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		48140 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		48141 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		48147 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		48156 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		48164 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		48180 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		48187 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		48199 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		48216 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		48218 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		48223 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		48224 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		48232 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		48238 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		48250 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		48251 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		48274 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		48282 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		48288 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		48312 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		48313 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		48315 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		48317 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		48321 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		48331 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		48335 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		48340 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		48347 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		48361 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		48365 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		48376 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		48379 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		48387 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		48410 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		48412 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		48414 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		48415 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		48421 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		48445 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		48451 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		48454 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		48464 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		48474 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		48476 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		48491 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		48498 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		48502 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		48509 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		48516 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		48519 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		48522 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		48527 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		48533 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		48542 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		48543 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		48550 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		48557 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		48570 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		48575 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		48578 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		48579 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		48581 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		48584 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		48585 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		48588 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		48615 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		48618 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		48635 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		48639 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		48644 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		48677 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		48680 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		48685 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		48687 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		48699 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		48701 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		48710 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		48714 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		48717 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		48726 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		48733 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		48737 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		48746 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		48753 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		48756 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		48759 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		48766 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		48769 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		48770 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		48775 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		48776 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		48789 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		48791 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		48800 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		48801 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		48830 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		48831 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		48832 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		48835 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		48848 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		48851 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		48866 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		48873 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		48878 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		48883 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		48888 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		48894 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		48900 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		48907 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		48908 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		48917 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		48922 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		48928 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		48940 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		48942 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		48947 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		48963 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		48990 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		48995 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		48996 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		48997 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		49002 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		49007 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		49024 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		49034 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		49037 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		49048 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		49055 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		49084 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		49094 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		49104 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		49109 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		49113 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		49115 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		49123 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		49125 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		49132 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		49133 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		49150 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		49182 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		49201 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		49209 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		49212 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		49234 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		49245 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		49248 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		49256 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		49259 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		49260 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		49263 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		49268 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		49275 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		49280 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		49281 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		49282 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		49290 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		49292 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		49295 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		49303 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		49305 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		49307 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		49319 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		49322 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		49325 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		49329 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		49331 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		49336 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		49338 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		49350 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		49351 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		49356 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		49386 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		49387 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		49419 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		49428 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		49459 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		49465 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		49476 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		49485 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		49495 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		49498 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		49505 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		49509 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		49524 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		49525 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		49532 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		49537 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		49545 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		49547 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		49548 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		49558 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		49578 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		49596 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		49599 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		49605 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		49606 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		49607 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		49609 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		49611 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		49613 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		49636 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		49637 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		49639 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		49647 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		49663 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		49666 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		49667 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		49673 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		49674 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		49676 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		49677 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		49678 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		49690 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		49701 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		49706 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		49723 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		49726 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		49733 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		49734 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		49735 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		49746 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		49747 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		49749 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		49761 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		49763 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		49785 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		49788 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		49790 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		49811 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		49812 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		49821 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		49825 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		49836 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		49841 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		49853 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		49854 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		49855 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		49861 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		49866 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		49884 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		49887 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		49890 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		49904 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		49910 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		49911 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		49916 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		49922 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		49924 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		49937 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		49941 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		49942 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		49953 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		49955 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		49957 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		49965 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		49972 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		49978 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		49979 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		49989 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		49995 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		50016 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		50027 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		50034 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		50037 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		50038 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		50039 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		50040 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		50043 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		50047 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		50051 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		50052 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		50057 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		50061 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		50063 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		50065 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		50081 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		50087 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		50095 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		50105 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		50132 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		50146 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		50152 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		50153 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		50156 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		50159 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		50177 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		50180 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		50186 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		50206 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		50210 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		50214 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		50234 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		50235 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		50244 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		50248 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		50251 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		50256 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		50259 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		50273 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		50276 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		50289 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		50292 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		50294 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		50306 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		50328 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		50329 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		50337 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		50338 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		50342 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		50345 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		50352 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		50361 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		50370 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		50371 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		50386 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		50395 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		50396 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		50397 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		50415 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		50423 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		50429 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		50438 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		50443 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		50453 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		50495 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		50510 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		50521 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		50531 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		50547 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		50549 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		50563 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		50571 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		50589 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		50603 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		50607 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		50610 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		50614 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		50644 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		50653 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		50678 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		50695 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		50718 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		50740 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		50747 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		50749 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		50753 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		50758 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		50766 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		50768 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		50777 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		50780 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		50785 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		50790 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		50805 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		50809 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		50814 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		50829 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		50830 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		50834 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		50837 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		50839 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		50841 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		50846 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		50848 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		50857 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		50859 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		50873 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		50877 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		50882 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		50884 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		50891 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		50895 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		50896 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		50900 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		50902 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		50910 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		50911 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		50919 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		50933 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		50935 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		50936 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		50952 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		50954 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		50960 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		50964 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		50965 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		50968 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		50974 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		50976 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		50978 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		50981 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		50982 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		50987 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		50989 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		50990 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		51002 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		51006 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		51010 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		51013 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		51015 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		51016 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		51024 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		51028 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		51030 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		51037 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		51040 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		51049 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		51076 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		51080 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		51082 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		51100 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		51109 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		51137 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		51142 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		51147 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		51149 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		51159 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		51170 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		51178 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		51183 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		51190 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		51196 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		51198 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		51200 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		51231 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		51240 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		51248 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		51249 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		51259 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		51263 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		51271 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		51285 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		51296 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		51297 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		51305 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		51319 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		51320 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		51324 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		51328 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		51347 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		51356 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		51370 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		51376 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		51382 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		51383 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		51385 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		51388 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		51390 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		51412 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		51414 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		51417 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		51430 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		51440 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		51442 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		51443 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		51445 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		51458 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		51466 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		51485 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		51491 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		51495 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		51510 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		51514 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		51517 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		51523 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		51534 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		51535 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		51536 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		51537 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		51541 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		51547 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		51555 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		51571 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		51575 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		51577 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		51587 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		51598 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		51602 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		51612 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		51644 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		51648 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		51661 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		51670 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		51682 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		51702 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		51703 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		51705 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		51720 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		51721 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		51728 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		51732 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		51735 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		51745 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		51749 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		51756 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		51758 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		51761 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		51772 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		51777 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		51783 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		51789 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		51790 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		51796 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		51803 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		51804 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		51805 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		51815 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		51816 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		51824 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		51835 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		51842 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		51844 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		51845 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		51849 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		51851 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		51854 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		51855 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		51868 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		51876 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		51883 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		51896 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		51903 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		51919 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		51923 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		51928 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		51961 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		51978 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		51980 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		51987 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		52009 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		52011 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		52013 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		52027 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		52047 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		52050 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		52057 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		52061 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		52062 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		52067 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		52071 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		52075 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		52078 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		52079 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		52083 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		52087 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		52098 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		52107 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		52119 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		52124 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		52136 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		52137 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		52146 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		52148 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		52151 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		52160 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		52162 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		52166 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		52181 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		52185 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		52191 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		52193 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		52202 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		52222 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		52224 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		52245 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		52249 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		52252 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		52253 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		52257 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		52260 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		52265 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		52272 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		52274 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		52279 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		52283 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		52296 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		52299 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		52304 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		52309 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		52316 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		52318 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		52324 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		52335 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		52337 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		52339 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		52340 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		52343 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		52344 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		52354 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		52358 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		52367 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		52372 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		52379 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		52395 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		52396 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		52398 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		52400 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		52407 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		52409 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		52410 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		52420 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		52423 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		52429 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		52435 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		52440 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		52457 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		52464 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		52471 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		52472 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		52480 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		52481 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		52485 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		52489 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		52491 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		52494 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		52500 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		52504 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		52514 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		52521 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		52527 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		52530 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		52533 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		52544 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		52547 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		52551 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		52553 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		52554 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		52557 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		52559 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		52561 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		52581 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		52586 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		52589 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		52592 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		52599 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		52603 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		52609 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		52620 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		52655 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		52669 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		52673 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		52675 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		52686 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		52692 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		52694 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		52701 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		52712 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		52720 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		52722 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		52727 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		52733 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		52738 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		52739 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		52740 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		52746 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		52756 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		52763 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		52765 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		52779 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		52780 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		52793 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		52817 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		52828 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		52853 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		52855 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		52867 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		52877 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		52921 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		52927 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		52928 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		52942 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		52944 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		52951 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		52958 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		52960 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		52975 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		52991 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		52998 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		53006 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		53009 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		53017 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		53055 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		53056 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		53066 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		53073 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		53078 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		53083 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		53084 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		53101 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		53103 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		53109 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		53111 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		53113 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		53121 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		53126 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		53129 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		53132 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		53138 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		53140 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		53151 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		53152 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		53154 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		53157 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		53172 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		53185 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		53186 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		53195 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		53200 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		53208 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		53217 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		53222 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		53224 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		53225 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		53228 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		53238 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		53243 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		53263 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		53264 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		53274 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		53275 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		53277 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		53285 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		53292 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		53293 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		53324 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		53327 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		53334 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		53336 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		53339 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		53347 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		53353 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		53355 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		53362 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		53363 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		53366 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		53373 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		53379 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		53384 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		53409 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		53410 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		53411 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		53419 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		53420 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		53453 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		53481 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		53516 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		53518 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		53521 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		53536 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		53541 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		53543 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		53551 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		53555 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		53558 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		53565 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		53569 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		53580 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		53596 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		53601 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		53642 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		53647 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		53650 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		53672 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		53684 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		53689 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		53690 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		53698 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		53705 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		53707 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		53718 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		53724 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		53728 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		53762 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		53766 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		53792 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		53802 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		53816 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		53843 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		53852 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		53857 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		53870 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		53871 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		53878 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		53879 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		53888 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		53894 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		53904 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		53907 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		53916 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		53932 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		53938 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		53940 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		53948 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		53960 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		53964 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		53968 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		53986 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		53990 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		54009 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		54011 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		54025 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		54029 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		54049 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		54055 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		54068 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		54071 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		54083 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		54084 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		54090 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		54091 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		54095 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		54099 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		54147 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		54154 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		54155 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		54163 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		54165 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		54166 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		54186 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		54188 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		54201 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		54225 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		54229 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		54231 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		54234 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		54251 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		54257 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		54281 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		54289 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		54290 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		54317 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		54344 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		54357 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		54360 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		54365 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		54369 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		54384 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		54388 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		54391 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		54395 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		54417 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		54418 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		54424 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		54439 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		54463 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		54467 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		54473 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		54478 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		54481 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		54485 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		54488 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		54493 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		54494 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		54496 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		54498 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		54510 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		54511 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		54515 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		54527 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		54550 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		54551 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		54563 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		54572 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		54574 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		54584 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		54597 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		54598 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		54604 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		54609 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		54622 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		54631 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		54632 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		54636 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		54637 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		54652 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		54654 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		54658 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		54661 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		54662 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		54682 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		54684 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		54688 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		54690 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		54691 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		54709 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		54719 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		54727 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		54732 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		54734 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		54737 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		54738 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		54765 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		54768 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		54781 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		54787 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		54792 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		54801 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		54806 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		54822 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		54828 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		54831 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		54835 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		54841 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		54848 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		54850 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		54852 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		54856 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		54867 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		54882 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		54887 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		54895 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		54897 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		54912 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		54919 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		54922 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		54926 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		54930 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		54934 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		54935 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		54942 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		54945 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		54946 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		54956 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		54960 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		54963 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		54967 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		54976 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		54987 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		54989 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		55000 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		55008 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		55029 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		55032 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		55049 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		55050 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		55053 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		55059 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		55062 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		55088 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		55090 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		55097 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		55118 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		55119 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		55129 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		55131 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		55146 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		55152 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		55160 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		55163 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		55166 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		55169 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		55171 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		55185 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		55193 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		55203 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		55209 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		55222 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		55225 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		55246 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		55256 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		55259 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		55279 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		55286 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		55290 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		55299 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		55300 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		55304 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		55305 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		55308 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		55316 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		55322 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		55323 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		55325 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		55335 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		55353 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		55354 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		55356 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		55364 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		55375 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		55376 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		55382 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		55391 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		55395 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		55411 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		55415 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		55416 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		55421 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		55423 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		55431 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		55433 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		55452 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		55454 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		55470 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		55479 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		55480 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		55481 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		55483 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		55500 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		55511 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		55532 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		55545 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		55550 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		55576 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		55577 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		55582 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		55588 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		55597 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		55599 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		55600 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		55628 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		55636 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		55637 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		55641 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		55644 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		55675 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		55679 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		55686 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		55692 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		55719 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		55740 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		55747 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		55757 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		55760 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		55765 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		55776 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		55793 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		55802 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		55803 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		55808 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		55823 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		55847 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		55850 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		55859 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		55870 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		55879 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		55883 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		55908 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		55916 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		55919 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		55934 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		55939 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		55944 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		55951 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		55963 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		55965 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		55976 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		55986 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		56005 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		56006 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		56014 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		56023 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		56033 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		56035 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		56039 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		56043 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		56061 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		56062 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		56072 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		56088 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		56089 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		56094 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		56103 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		56108 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		56111 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		56119 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		56123 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		56137 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		56143 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		56145 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		56146 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		56150 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		56152 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		56156 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		56158 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		56172 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		56185 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		56186 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		56188 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		56191 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		56195 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		56198 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		56203 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		56229 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		56232 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		56234 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		56237 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		56250 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		56258 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		56267 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		56271 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		56272 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		56278 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		56279 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		56283 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		56289 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		56291 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		56293 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		56296 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		56297 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		56300 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		56309 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		56310 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		56324 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		56328 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		56330 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		56333 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		56342 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		56357 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		56361 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		56364 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		56368 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		56372 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		56374 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		56386 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		56388 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		56391 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		56392 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		56401 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		56410 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		56413 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		56414 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		56416 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		56427 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		56441 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		56446 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		56468 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		56479 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		56485 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		56492 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		56504 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		56510 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		56513 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		56519 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		56525 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		56533 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		56536 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		56562 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		56563 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		56564 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		56566 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		56567 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		56574 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		56575 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		56576 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		56586 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		56588 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		56591 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		56602 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		56611 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		56613 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		56625 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		56627 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		56629 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		56649 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		56669 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		56670 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		56672 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		56677 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		56682 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		56688 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		56693 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		56694 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		56703 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		56709 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		56710 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		56718 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		56725 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		56733 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		56745 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		56747 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		56750 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		56759 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		56771 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		56778 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		56779 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		56781 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		56782 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		56783 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		56792 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		56797 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		56798 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		56801 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		56802 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		56810 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		56816 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		56830 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		56831 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		56833 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		56848 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		56865 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		56869 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		56882 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		56884 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		56888 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		56890 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		56891 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		56892 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		56897 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		56900 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		56902 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		56910 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		56921 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		56928 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		56933 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		56946 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		56976 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		56980 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		57000 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		57005 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		57009 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		57017 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		57019 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		57020 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		57026 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		57032 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		57034 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		57037 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		57044 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		57048 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		57051 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		57052 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		57057 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		57066 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		57071 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		57080 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		57093 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		57097 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		57098 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		57105 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		57107 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		57113 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		57119 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		57120 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		57123 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		57129 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		57133 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		57143 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		57151 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		57169 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		57171 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		57175 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		57193 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		57204 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		57206 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		57212 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		57239 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		57240 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		57248 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		57252 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		57261 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		57262 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		57263 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		57264 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		57265 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		57274 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		57277 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		57285 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		57298 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		57300 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		57339 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		57343 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		57345 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		57347 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		57349 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		57357 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		57371 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		57376 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		57392 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		57394 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		57406 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		57413 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		57416 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		57421 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		57426 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		57431 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		57435 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		57443 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		57446 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		57460 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		57463 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		57471 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		57473 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		57477 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		57485 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		57490 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		57496 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		57501 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		57508 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		57515 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		57523 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		57539 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		57545 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		57551 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		57555 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		57556 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		57572 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		57577 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		57581 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		57586 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		57587 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		57588 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		57600 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		57605 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		57640 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		57646 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		57650 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		57654 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		57665 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		57669 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		57675 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		57716 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		57718 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		57719 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		57720 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		57731 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		57744 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		57759 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		57766 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		57790 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		57792 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		57809 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		57812 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		57816 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		57817 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		57819 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		57822 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		57827 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		57834 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		57837 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		57849 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		57861 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		57873 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		57891 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		57892 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		57893 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		57894 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		57895 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		57896 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		57916 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		57923 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		57927 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		57931 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		57936 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		57949 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		57950 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		57952 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		57979 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		57986 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		57988 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		58002 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		58005 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		58017 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		58031 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		58035 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		58048 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		58050 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		58084 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		58085 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		58090 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		58092 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		58093 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		58094 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		58098 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		58101 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		58109 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		58131 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		58137 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		58143 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		58172 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		58180 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		58186 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		58195 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		58207 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		58212 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		58214 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		58220 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		58223 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		58241 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		58242 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		58243 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		58250 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		58251 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		58255 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		58257 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		58260 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		58267 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		58271 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		58273 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		58284 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		58299 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		58300 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		58311 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		58326 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		58328 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		58335 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		58354 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		58358 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		58370 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		58374 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		58384 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		58400 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		58402 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		58404 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		58408 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		58409 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		58411 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		58419 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		58423 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		58424 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		58428 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		58438 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		58442 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		58456 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		58462 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		58472 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		58480 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		58504 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		58506 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		58509 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		58514 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		58516 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		58518 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		58530 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		58535 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		58541 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		58558 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		58561 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		58565 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		58590 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		58592 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		58595 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		58598 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		58604 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		58610 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		58620 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		58638 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		58645 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		58647 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		58654 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		58657 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		58659 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		58668 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		58679 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		58680 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		58694 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		58702 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		58704 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		58725 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		58734 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		58751 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		58755 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		58760 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		58762 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		58775 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		58776 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		58798 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		58804 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		58807 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		58809 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		58811 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		58818 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		58822 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		58828 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		58842 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		58844 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		58846 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		58848 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		58854 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		58872 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		58874 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		58885 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		58886 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		58893 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		58899 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		58901 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		58929 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		58931 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		58936 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		58944 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		58948 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		58952 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		58957 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		58958 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		58960 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		58965 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		58982 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		58993 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		58997 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		59009 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		59013 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		59016 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		59019 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		59036 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		59049 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		59058 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		59068 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		59073 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		59075 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		59082 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		59083 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		59087 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		59090 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		59095 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		59102 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		59109 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		59118 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		59126 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		59137 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		59141 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		59144 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		59147 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		59150 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		59171 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		59174 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		59187 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		59190 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		59192 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		59198 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		59202 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		59206 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		59215 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		59220 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		59222 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		59239 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		59241 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		59244 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		59249 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		59252 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		59264 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		59277 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		59279 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		59280 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		59291 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		59298 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		59301 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		59306 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		59308 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		59317 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		59319 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		59344 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		59346 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		59347 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		59348 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		59352 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		59354 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		59360 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		59376 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		59378 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		59384 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		59385 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		59392 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		59404 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		59406 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		59421 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		59428 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		59434 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		59435 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		59443 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		59464 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		59466 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		59471 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		59477 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		59489 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		59496 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		59501 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		59505 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		59515 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		59545 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		59563 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		59570 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		59594 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		59607 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		59620 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		59626 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		59627 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		59632 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		59638 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		59639 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		59646 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		59657 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		59661 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		59687 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		59688 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		59710 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		59711 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		59714 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		59717 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		59722 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		59733 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		59735 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		59748 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		59750 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		59752 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		59754 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		59758 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		59762 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		59773 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		59780 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		59781 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		59787 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		59791 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		59798 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		59802 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		59804 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		59813 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		59826 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		59841 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		59845 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		59849 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		59853 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		59855 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		59856 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		59867 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		59871 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		59873 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		59879 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		59883 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		59884 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		59887 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		59890 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		59895 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		59898 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		59902 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		59905 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		59911 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		59919 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		59925 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		59927 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		59928 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		59929 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		59944 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		59948 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		59959 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		59966 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		59973 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		59976 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		59984 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		59986 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		59988 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		60001 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		60010 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		60015 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		60027 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		60032 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		60039 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		60052 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		60056 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		60060 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		60061 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		60065 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		60074 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		60092 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		60095 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		60104 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		60110 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		60111 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		60115 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		60121 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		60122 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		60132 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		60133 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		60139 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		60140 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		60147 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		60164 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		60168 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		60170 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		60172 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		60183 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		60185 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		60187 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		60188 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		60197 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		60204 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		60205 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		60210 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		60211 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		60217 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		60220 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		60224 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		60228 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		60235 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		60251 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		60252 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		60253 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		60256 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		60259 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		60269 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		60286 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		60290 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		60292 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		60300 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		60307 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		60309 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		60310 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		60311 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		60314 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		60322 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		60335 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		60341 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		60348 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		60351 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		60366 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		60367 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		60368 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		60378 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		60382 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		60386 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		60392 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		60399 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		60407 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		60409 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		60414 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		60427 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		60429 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		60433 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		60438 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		60451 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		60456 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		60459 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		60460 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		60473 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		60484 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		60487 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		60490 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		60491 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		60493 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		60495 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		60500 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		60507 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		60510 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		60512 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		60516 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		60518 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		60522 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		60523 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		60533 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		60534 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		60535 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		60536 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		60543 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		60570 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		60579 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		60591 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		60592 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		60610 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		60628 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		60650 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		60656 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		60659 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		60667 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		60679 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		60681 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		60694 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		60696 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		60698 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		60703 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		60706 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		60707 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		60709 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		60713 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		60717 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		60730 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		60777 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		60791 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		60797 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		60800 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		60810 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		60817 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		60827 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		60835 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		60844 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		60854 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		60859 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		60864 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		60897 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		60903 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		60905 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		60915 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		60920 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		60922 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		60924 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		60946 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		60950 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		60956 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		60963 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		60965 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		60966 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		60977 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		60981 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		60988 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		60996 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		61000 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		61003 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		61011 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		61019 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		61023 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		61038 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		61040 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		61045 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		61049 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		61055 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		61056 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		61057 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		61059 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		61064 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		61073 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		61079 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		61088 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		61089 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		61092 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		61094 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		61103 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		61106 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		61108 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		61119 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		61122 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		61123 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		61125 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		61127 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		61134 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		61135 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		61141 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		61153 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		61160 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		61162 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		61166 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		61168 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		61172 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		61183 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		61191 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		61192 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		61193 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		61196 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		61209 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		61217 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		61219 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		61222 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		61227 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		61236 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		61240 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		61242 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		61247 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		61251 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		61264 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		61286 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		61301 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		61302 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		61326 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		61329 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		61332 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		61333 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		61341 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		61355 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		61358 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		61380 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		61386 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		61411 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		61419 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		61420 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		61427 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		61429 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		61439 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		61441 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		61445 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		61452 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		61456 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		61492 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		61496 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		61522 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		61528 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		61542 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		61544 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		61546 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		61547 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		61571 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		61575 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		61589 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		61599 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		61600 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		61601 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		61608 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		61610 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		61615 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		61618 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		61620 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		61623 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		61627 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		61634 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		61638 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		61641 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		61645 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		61658 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		61683 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		61687 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		61688 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		61691 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		61693 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		61703 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		61716 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		61720 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		61727 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		61736 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		61739 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		61746 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		61748 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		61749 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		61752 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		61753 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		61761 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		61767 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		61768 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		61785 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		61790 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		61803 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		61818 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		61825 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		61829 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		61836 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		61842 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		61843 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		61851 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		61856 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		61858 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		61873 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		61875 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		61877 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		61893 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		61914 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		61925 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		61948 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		61952 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		61954 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		61955 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		61966 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		61974 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		61988 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		61992 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		61995 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		61996 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		62002 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		62005 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		62006 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		62008 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		62019 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		62035 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		62036 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		62040 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		62047 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		62048 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		62054 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		62086 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		62103 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		62105 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		62109 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		62119 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		62124 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		62125 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		62142 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		62150 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		62151 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		62152 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		62153 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		62161 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		62183 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		62184 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		62185 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		62195 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		62198 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		62199 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		62204 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		62210 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		62220 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		62235 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		62241 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		62252 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		62259 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		62262 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		62265 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		62270 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		62276 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		62277 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		62278 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		62286 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		62292 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		62310 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		62315 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		62319 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		62333 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		62334 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		62344 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		62351 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		62353 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		62354 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		62356 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		62366 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		62376 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		62380 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		62406 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		62413 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		62423 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		62432 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		62442 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		62443 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		62444 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		62445 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		62447 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		62451 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		62454 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		62457 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		62463 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		62480 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		62484 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		62490 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		62505 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		62506 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		62507 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		62510 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		62526 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		62540 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		62546 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		62549 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		62568 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		62598 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		62612 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		62615 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		62617 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		62623 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		62625 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		62626 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		62629 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		62637 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		62638 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		62640 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		62641 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		62645 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		62657 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		62660 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		62664 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		62667 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		62671 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		62680 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		62685 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		62688 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		62689 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		62691 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		62701 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		62709 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		62718 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		62719 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		62737 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		62751 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		62753 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		62755 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		62759 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		62760 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		62761 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		62763 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		62764 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		62767 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		62770 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		62794 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		62799 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		62806 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		62812 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		62816 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		62818 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		62838 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		62842 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		62847 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		62855 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		62877 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		62881 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		62890 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		62892 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		62899 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		62915 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		62919 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		62921 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		62923 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		62936 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		62937 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		62940 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		62960 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		62964 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		62968 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		62981 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		62982 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		62986 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		62991 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		62994 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		62999 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		63002 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		63003 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		63008 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		63012 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		63018 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		63024 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		63033 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		63036 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		63044 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		63052 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		63061 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		63064 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		63091 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		63097 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		63101 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		63107 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		63114 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		63117 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		63121 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		63159 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		63162 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		63170 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		63178 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		63183 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		63184 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		63203 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		63206 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		63207 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		63212 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		63236 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		63240 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		63251 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		63266 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		63269 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		63286 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		63309 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		63311 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		63312 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		63315 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		63322 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		63335 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		63346 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		63349 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		63351 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		63353 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		63357 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		63370 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		63381 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		63399 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		63417 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		63422 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		63423 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		63436 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		63441 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		63448 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		63452 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		63466 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		63468 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		63473 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		63487 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		63494 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		63497 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		63507 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		63509 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		63514 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		63516 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		63522 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		63526 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		63555 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		63561 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		63567 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		63569 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		63572 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		63591 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		63598 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		63599 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		63601 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		63610 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		63611 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		63619 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		63629 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		63644 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		63655 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		63670 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		63674 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		63675 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		63679 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		63680 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		63691 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		63700 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		63703 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		63708 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		63715 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		63730 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		63733 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		63734 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		63740 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		63741 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		63743 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		63748 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		63753 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		63758 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		63760 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		63778 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		63784 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		63794 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		63799 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		63814 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		63820 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		63846 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		63851 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		63861 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		63865 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		63869 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		63872 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		63882 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		63883 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		63885 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		63893 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		63897 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		63904 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		63910 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		63924 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		63926 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		63935 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		63942 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		63943 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		63944 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		63954 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		63963 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		63971 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		63974 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		63990 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		63996 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		63999 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		64006 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		64007 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		64008 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		64009 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		64010 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		64022 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		64034 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		64035 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		64084 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		64095 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		64096 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		64100 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		64110 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		64111 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		64143 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		64146 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		64148 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		64151 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		64168 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		64171 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		64182 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		64224 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		64239 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		64241 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		64244 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		64248 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		64250 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		64263 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		64274 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		64275 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		64279 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		64282 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		64290 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		64293 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		64296 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		64298 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		64299 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		64304 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		64316 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		64319 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		64322 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		64333 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		64342 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		64343 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		64346 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		64348 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		64354 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		64356 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		64361 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		64364 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		64367 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		64387 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		64392 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		64394 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		64396 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		64400 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		64405 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		64410 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		64413 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		64417 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		64424 => STD_LOGIC_VECTOR(to_unsigned(43,8)),
		64439 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		64448 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		64456 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		64457 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		64462 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		64480 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		64493 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		64496 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		64497 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		64499 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		64500 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		64501 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		64508 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		64509 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		64513 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		64522 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		64523 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		64539 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		64540 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		64542 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		64548 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		64565 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		64566 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		64572 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		64574 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		64584 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		64599 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		64603 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		64604 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		64611 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		64612 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		64617 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		64620 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		64621 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		64625 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		64640 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		64645 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		64659 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		64660 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		64667 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		64669 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		64685 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		64695 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		64698 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		64701 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		64707 => STD_LOGIC_VECTOR(to_unsigned(108,8)),
		64709 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		64718 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		64730 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		64733 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		64737 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		64744 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		64773 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		64774 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		64776 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		64779 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		64799 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		64808 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		64834 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		64839 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		64846 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		64848 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		64853 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		64877 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		64890 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		64897 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		64904 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		64909 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		64916 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		64917 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		64919 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		64928 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		64930 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		64931 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		64943 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		64945 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		64947 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		64950 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		64954 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		64955 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		64963 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		64975 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		64982 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		64983 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		64989 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		64990 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		64991 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		65018 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		65022 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		65023 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		65034 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		65036 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		65039 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		65045 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		65054 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		65055 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		65056 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		65065 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		65071 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		65081 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		65085 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		65088 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		65094 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		65098 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		65101 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		65110 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		65151 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		65161 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		65163 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		65164 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		65180 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		65187 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		65189 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		65194 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		65212 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		65219 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		65221 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		65227 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		65236 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		65256 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		65260 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		65264 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		65274 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		65286 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		65292 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		65308 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		65309 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		65316 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		65317 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		65320 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		65326 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		65327 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		65329 => STD_LOGIC_VECTOR(to_unsigned(62,8)),
		65354 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		65365 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		65372 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		65384 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		65403 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		65409 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		65412 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		65414 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		65423 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		65430 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		65434 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		65439 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		65452 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		65472 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		65479 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		65488 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		65491 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		65505 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		65508 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		65519 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		others => (others => '0')
	);

	COMPONENT project_reti_logiche IS
		PORT (
			i_clk : IN STD_LOGIC;
			i_rst : IN STD_LOGIC;
			i_start : IN STD_LOGIC;
			i_w : IN STD_LOGIC;

			o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_done : OUT STD_LOGIC;

			o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_mem_we : OUT STD_LOGIC;
			o_mem_en : OUT STD_LOGIC
		);
	END COMPONENT project_reti_logiche;

BEGIN
	UUT : project_reti_logiche
	PORT MAP(
		i_clk => tb_clk,
		i_start => tb_start,
		i_rst => tb_rst,
		i_w => tb_w,

		o_z0 => tb_z0,
		o_z1 => tb_z1,
		o_z2 => tb_z2,
		o_z3 => tb_z3,
		o_done => tb_done,

		o_mem_addr => mem_address,
		o_mem_en => enable_wire,
		o_mem_we => mem_we,
		i_mem_data => mem_o_data
	);


	-- Process for the clock generation
	CLK_GEN : PROCESS IS
	BEGIN
		WAIT FOR CLOCK_PERIOD/2;
		tb_clk <= NOT tb_clk;
	END PROCESS CLK_GEN;


	-- Process related to the memory
	MEM : PROCESS (tb_clk)
	BEGIN
		IF tb_clk'event AND tb_clk = '1' THEN
			IF enable_wire = '1' THEN
				IF mem_we = '1' THEN
					RAM(conv_integer(mem_address)) <= mem_i_data;
					mem_o_data <= mem_i_data AFTER 1 ns;
				ELSE
					mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns;
				END IF;
			END IF;
		END IF;
	END PROCESS;

	-- This process provides the correct scenario on the signal controlled by the TB
	createScenario : PROCESS (tb_clk)
	BEGIN
		IF tb_clk'event AND tb_clk = '0' THEN
			tb_rst <= scenario_rst(0);
			tb_w <= scenario_w(0);
			tb_start <= scenario_start(0);
			scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
			scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
			scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
		END IF;
	END PROCESS;

	-- Process without sensitivity list designed to test the actual component.
	testRoutine : PROCESS IS
	BEGIN
		FOR i IN 0 TO N_EVENTS - 1 LOOP
			mem_i_data <= "00000000";
			IF do_reset(i) = '1' THEN
				WAIT UNTIL tb_rst = '1';
				WAIT UNTIL tb_rst = '0';
				ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure;
				ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure;
				ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
				ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
				ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset done != 0 )" severity failure;
				ASSERT enable_wire = '0' REPORT "TEST FALLITO (postreset enable_wire != 0 )" severity warning;
				ASSERT mem_we = '0' REPORT "(mem_we != 0 )" severity failure;
			END IF;

			WAIT UNTIL tb_start = '1';
			ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure;
			ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure;
			ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
			ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure;
			ASSERT tb_done = '0' REPORT "TEST FALLITO (poststart done != 0 )" severity failure;
			ASSERT enable_wire = '0' REPORT "TEST FALLITO (poststart enable_wire != 0 )" severity warning;
			ASSERT mem_we = '0' REPORT "(mem_we != 0 )" severity failure;
			WAIT UNTIL tb_done = '1';
			--WAIT UNTIL rising_edge(tb_clk);
			WAIT FOR CLOCK_PERIOD/2;
			ASSERT tb_z0 = std_logic_vector(to_unsigned(registers_check(i, 0), 8))	REPORT "TEST FALLITO (Z0 ---) found " & integer'image(to_integer(unsigned(tb_z0))) & " Expected " & integer'image(registers_check(i, 0)) severity failure;
			ASSERT tb_z1 = std_logic_vector(to_unsigned(registers_check(i, 1), 8))	REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z1))) & " Expected " & integer'image(registers_check(i, 1)) severity failure;
			ASSERT tb_z2 = std_logic_vector(to_unsigned(registers_check(i, 2), 8))	REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z2))) & " Expected " & integer'image(registers_check(i, 2)) severity failure;
			ASSERT tb_z3 = std_logic_vector(to_unsigned(registers_check(i, 3), 8))	REPORT "TEST FALLITO (Z3 ---) found " & integer'image(to_integer(unsigned(tb_z3))) & " Expected " & integer'image(registers_check(i, 3)) severity failure;
			ASSERT tb_done = '1' REPORT "TEST FALLITO (done = 0 )" severity failure;
			WAIT FOR CLOCK_PERIOD/2 + 10 ns;
			ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure;
			ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure;
			ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
			ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure;
			ASSERT tb_done = '0' REPORT "TEST FALLITO (postdone done != 0 )" severity failure;
			ASSERT enable_wire = '0' REPORT "(postdone enable_wire != 0 )" severity warning;
			ASSERT mem_we = '0' REPORT "TEST FALLITO (mem_we != 0 )" severity failure;
		END LOOP;
		wait FOR CLOCK_PERIOD * 2;
		REPORT "SUCCESS";
		finish;
	END PROCESS testRoutine;

END randomtb;

