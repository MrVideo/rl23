
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;
USE std.env.finish;

ENTITY random_tb IS
END random_tb;

ARCHITECTURE randomtb OF random_tb IS
	CONSTANT CLOCK_PERIOD : TIME := 100 ns;
	SIGNAL tb_done : STD_LOGIC;
	SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
	SIGNAL tb_rst : STD_LOGIC := '0';
	SIGNAL tb_start : STD_LOGIC := '0';
	SIGNAL tb_clk : STD_LOGIC := '0';
	SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL enable_wire : STD_LOGIC;
	SIGNAL mem_we : STD_LOGIC;
	SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL tb_w : STD_LOGIC;

	CONSTANT SCENARIOLENGTH : INTEGER := 40549;
	CONSTANT N_EVENTS : INTEGER := 1000;
	SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)		:= "0100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)	:= "0100011111111111111111100000000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000001111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000010000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000100011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000001111111111111110000000000000000000001111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000001111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000001000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000001000111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111100000000000000000000000111111111111111110000000000000000000000011111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000001111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111111000000000000000000001000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000001111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000010111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100011111111111111111000000000000000000000000111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000001111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000010001111111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000001111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000000001111111111111111110000000000000000000010000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000000111111111111111110000000000000000000000001111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111100000000000000000000100000111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000001111111111111111000000000000000000000000011111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000001111111111111111000000000000000000001011111111111111111100000000000000000000011111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000011111111111111110000000000000000000000011111111111111110000000000000000000000011111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000001111111111111111000000000000000000001011111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000001111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000101111111111111111110000000000000000000000001111111111111111110000000000000000000010001111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000010011111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000001001111111111111111000000000000000000000001111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111100000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000001000011111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000001111111111111111100000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111100000000000000000000100001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000000111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000010011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000010001111111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111000000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000001111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000101111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111100000000000000000000011111111111111100000000000000000000000111111111111111111000000000000000000001000011111111111111110000000000000000000000001111111111111111110000000000000000000000111111111111111110000000000000000000000011111111111111110000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000100001111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000100000111111111111111111000000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000100000111111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000001111111111111111110000000000000000000010011111111111111111100000000000000000000000001111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000011111111111111111100000000000000000000100011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000111111111111000000000000000000000111111111111111110000000000000000000000000111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111110000000000000000000000111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000100111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000001001111111111111111110000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111000000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000011111111111111110000000000000000000001111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000011111111111111111100000000000000000000000001111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000001111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111000000000000000000000000111111111111111110000000000000000000010111111111111111110000000000000000000000000111111111111111100000000000000000000000011111111111111111100000000000000000000100001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000011111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000011111111111111111100000000000000000000";
	SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)		:= "0100001010011001111010111110000001001011011001110010110011011010111100101110001011011000110110000011000010000000101011101101010100110001101101100110101110001000011100010111110101010111111011011110101111110100101011000101010001100100110110001000010011010111100001010101100100111101111111001011101111010110101101000011101111000101100110111100100111011101111100011011100010010001101111100111010100001010100001011010010101001011100111100001010000100001100010111000111110101110101100110110110001100101101101011001100011111000000010100001001100100111011101110000111010010010000001101000100000001110100110110100101111011111001100010111110001110001101000101101010011011001011110000110010010110000001000001101010000101100100011000001101001001101011000010000101100000010100010000111000001110010001011101100010010001000111010111001100110101001001010001101001110111011111000101101111011100101100111101101011010001101010011101110011010100101011010110010001111100011000001100001101011111001011101000001011000111001000001010011011101001001011000110010011111000110101101011100011010100010101011111010001010100011111011011010111011100011010100010011110111101001010111110110101111000011000110100111001101011110101010010100111110011010010111101110111111110010000101001000101101101100101111001101001000010111110101111101001001011000111101011110010001010111000110000111111111101111100100001110101010110000001110011110111010111000111111011110010011010100010111110010110101111011001101111100100100010101001101011100010111111100001000000110010000010010011100010111010001110100110011011110000101111100100100011011010001110100010010000011011011010100100000100100110100110111100001001010100011001000000000100010010000010101101100010110000011110100011101111110001111010011001101010011011111011011111110110111111101110111110001010110100011111001111101010100001000100100101001010111000010111110110010111000100100111011000101001111100111001111010110111101000001000111001001010111010100111000110110101000100000101101100010110010001110011010110001010011001111011101101010011011010010100001001001000000100101001110101101111101010101010110101011000101110111100111011111101000101110111010111000001101010110011110101001000010101111110101110111100100111000110110010000110000101111100000001001010110001100010110010011100010010110111010000011000111110111001000011110101000001101011011011110011110101110011000110010101010101100111101001001100001001110111011111010111110101001010010100111011011110111110010101100100101000010010000011100110100000111111010100100001110000001010111000011100111111010101001100010000100100000111110010101110011110011100011100010011101010000010100111111001110000100100010000110000010010000010101000010011110111001001111101110011110011011000011111111111111011000010100000101010011010100100111011101001110010000101001000010110101101111101011110010100000001110011110001101010101100101000011100111011111111011110001111000010011000111110001000000001100000001000100110011101110110000110000011001000100011110111001111100011101101100101011110010100000111010101010011100001100000111110110101000100100101010111110110110001000011101100100000001110011011001010011010011010000111110011111110010100111001001000010011000001101100100101010001111010001010100001101001010001111110011010100101001001100110111100000000100101101001000000110001101001111111110000110000000100100110100100101000000010001110110011101100011110000101110001101011011101110111110100010110101111010100010000011111101000110111010110010110011101011110011010010011110010101111110011100011100101001100101110000111101011000000010101111011110111000110111010010001011001101011101001110001000100000011011101010010010101010101110111001001000011000110001100101000001111001110011010111101101111111100010000101101111011001011011000000100101111000100011101000100011111111001101111010111110010011110011100010111111010010000001110010010111011001110001001000011000011100110100011111010100001100000111000110111101101011111000001100100001110111011110110101000000111010011000101110000000010110011100001001001011100111011110000001101010101010100101000000111010101101001111011110100010101001110110011111110001011110101111000101100110111001000010000010001010010000011100010110010000101000001001100011000001100011010010010101100100100001110011011111000111111001010100100011001110101111010000011101001010010111001010111010010110100000111011111101010101111100011101011110001100100000100001100110110100110111111100011101111110010011000000000010100000010010000111101100111100010100010100001010011110100000000101011110110111001001111010110101000011001000101111011101110000101101101010001011001100110001101101001001110100001011010010100100011001100110000100001110100101111010000100111011111110010001101011111011011110010000000011010110000101000011011000010011110100011111010101010101100110101010101001000000000010000110111001001010011110011110111101110101010010110100110101101011010111001010101100111000100100001100010101100000010100110000001000110101110010011110100111010010001101100110111111100000001000010100010010011101111011110110001000000110110011111101010010010110001111010001000100101000111010111111101010000110000010101111101100100011111011011001111111100001011101100010001101111100100010001011010111011101010110010101011101101010001110111101011110101101010100000111110101001100111011011111011010111011110110101001101001100100001000101111110100111100100111010011111101110011101010110000101100111101110001000010000000010100011100110010110011100111001101111010100111000101010100011100110101011110011111100101001010001111000111010000000010000110000110111010001100010001110101010000011100110000100111100110000100110100000001101011001010010001111001100100000001000000100110000001011110101001110011110001100010100011000101000000011101001011010011101010110100001000111101000101011110100011010101111010010000100110101100110111011111010010101001001011011000111000010010001100001000101011101000010000001101011110110110111110110110100110000000000011100011011001011001011001100101010111010101011000111110111011111110000110000100001010010111110000111001110110111000100010101101001110001000010010001010110011100110101111010010011000001000111110100000001010101111110110010010010011001001001101000000110000101110100001000100010111111111001011101111110100111000100000111011101010100100000100100101101100110111001111000110111010001000000100011010001110100111000111000101000110101100001100000111100001000110111000111001100001110000101101001111101101010001010111110110101010001011111011101110011100111110010000111011001000100100011110101111011111001100011011001011101011011111100000111110101111111101000001000101100111011010001100010001111010000100000000101000000011010110111110100011101001010100011110100100010000001100000000100111111100010001010111111011001010011010101101110101110011100011011010100110010100100000100001001111111101110011001010111000111101000111010111000110100111011100101011110110100001111110101000001001011110001011110000010101010010111001100011100001001011000010010011011011011101110111000110101101010000010001100010101011111110101100111000011010101100011000111110011111011100111000001001000100010101100110011010011011110010011100110001100000110001000111111100110001000010111001000011011001010100000001011000111101101111100110100011000011111110011111011111001111100011111001001110100011010110010010100101010010000111101010001011100100101000110010100000101110100001111000100110110001000011001110100110110110011001010001101110110010101000111100000110101001011100101010110101110001000111011000101101110100001110100010101110001000101001101100000000010000000110110111001001111010001111101010001101110011111000111110011011110101101100111010001101001000111010001101000110000101100110010101101110000010011101011011011001101010100011101101100011110010011001000010010110100001101100010101100110011000011110010011001100100101001110001011000110000111001011011011100111101101110101000100000001011100111011111001011101001001010011010110011111101101100111100110111100011100100101111001001010011100001000010001100000000111110010101101100001001000001010110000100001011101011101101000010000110010101100001010111101010110110001101001000111000101010101101110001000100001101110011100100101011001000111110010001101000001111100111001101001101011000001000011000010001110101110100101100010100100100100111011100000100011000001100100010101100111000100111111101111100011110000110011011110101000110111011111110000010110001101110000100100000011011111010101101111110110011111001000110101101111001100001100111110101101010000011000100100010000011011011101110011011111010110011011111110001100011101111100110000110000111110100111100011110000001001001001110001000010100100011000000100110011000101000000111000001011111011111010101011111111101100001001100100101010111111100011100110010011010011011001100111010110111010100011100010011101101000010010010011001111100001001111110101111000010001111000111011101101110010010010010011010001010110100111110000110011000101000001110110110101110110010001001011011000111110101010011110100101100100111101101100100111001010001110000010110111100010001110010101101111101111010011101111110011010011010111101111100010110001000101111101101101100010110100111011111010110111001011010010100001001010000101001011001110100011011011011000111101010101000110000111110011011100010000001010100001101111111101010100010010100101101101111101100000010010101011011100101101100011101001101110111000101100000010001011011101000111100110101110110111001111100100001010110000001110101001000111111001110111111110011101111111010010111000011111011111101010010100010011101101111000111010001010001000001000000110000010001101100111111110101001101011001110111111010100001100000110010111011100001100001110110100011101001110011110101110001011001011010111000001100100101111110100011100010100011011011000010011010100010000011010100111000110010111010110010111110010111101010110101000001100110001001100000010110011111111010011101111111100111101011110101101010000011110111010110010001000111101111000100010000001111111100011110010011001100011000111110011111101010110000010101111110101111101111111010000001011100111111000111010111111101000101111001001010000001000111001001011110101011111110000101001111000101101001010001010001101011001010010011011011001101111111010011010101010101110011000110101111111011110101110001100100110011101110110010110010010011001000000111111000010101101111001100101101110001001001100010000011111000000000111010110110000110010101101001101101000001000101101001001010111010011000110100101001000100010100101001101101101010110110111101000011110110110100001110100111111011111101100101110010100100001100001110010100001011000100111111101110010100000001100001001100001110011100100100111000110011001101101111011101001110100001100100000000010001010100110010001001001000001010110000011101110100101011011100101011101010110100111101011100110111110101001110000000011101011010110111111111111101010100111101100110110000001100010110111100101100011001011011101100011011000010001100011101100100001000001101010000100100110000110100101111001100001110000011011100011000110001010010111000000110001011001100000000111011001110110111011110101110001011000111100000111000000100010001011110100101100100000000110111110110110010010001101111000110100110110011010101100100010101111101010100011010010000101000010111010111111001111010011100100001100000110110101100011011000010111010110101111100011010000110010010101111011010000101010011011100110011001001011101100000110101011010111000001010101111101000100010010100100100001100000010111010111100100110001010001110011000001110000000101101110001011011011010001010000000110101110101011110110011010001010011001111111110011011101111010000110110011100000010111110110110111110110010111111101011011001111000101111011111111101010110001101100000001011110100100101001011111110110110110110100111010101101010001011101111000001111101010111001111110100111000001110110011111010110100011100111100101011100011010111011101011001010110011100010011111111111110101110101011011000010001011000100101011011010011100111111110011001001010111011010101111110110010110001010011101000011011011011001110101111011101010001111101010101000101001101111000101010001110100000100010000011100101001100110010011000100011000111110101011010100111010011111110110101110101101011010101111010101110101010011101010000111011000001110010101101110001110010011100010111101111101100011111011000110110011011100100110001101000001010110001011001011111010001010010101110100000010010001001011000110000010110011000001110000110101010110010111001111111111100010100011101000011001001111001110111101000011110001010100100011111101101000011000111101011101010011111110101101100100000110010011111001001101010000110000011010111101111001011111100011110000111111110100000111001010001010000011101101111011001000010110011001110011110110101011101000011000011101000111111111001101001001111000110110101010101101000110000111001110010101101010101111111010011110101101001001000100011101111011111111101011101110000111100101101011001110111001111010111001011010011000001010101010001100001011110010010100010010001110101100011010110110110100011000111100101110111100001110000110010101011010100011011011011101111010110100100110001111110011000110101100010100110011101101011110111100101001011100000111101001101110101000111110101110100101000110011110000111101100011001100001000011010011010010101100000010011111000010110101000101010000110110000011110110001001111101110100101000101010100101010011011000101010111010111010001100001001011011000010100001100100110010000010001010011000110111000111011001110111011101111110100100000010100011111111100111111001101100101011011111011100110100110110110110010000110010001110100010100101010111111101110110010101001011001101000000111000111100011101100101011110101100011000000111111101110110000001101010110010111010011111000011110010111010111110110110001100001000010000001001100010101001110100010001110001011100011100101001010011011000110010010100100001001001101100101001000010011010101110111101111111001000010011011001111011100001110100110011010111100001110100101111111011010000100000100101111010001010010100111110100101001111001011110100110000100011011110100000110100111011001100001111110101100110000000010101010000000011001100000111100010101111100000000010001111000100010010000101001011011100000011011001100100010111100101001100100111000111101101011000111010001011011100100110101001000000110001100110000011011010101111011100100010101111110110010000111000010010001010010001101010000010000010111110000100011101001010001010001001110110000000101111011000001101100010101101001000111010010100011001010111110101011101101001011110101011111101100100001011010010110110101001111010000010110101101111101001010010100100101001110001110001000011100111100000011010011101000011010000001010001010100110010110011010100100111100111110100001110001101101001111100101110001100100101000111100111010100111000110110000111010110101111111100001000100001000010101001000101100010011000111000010000110001010001101010011000111110111011111011000010110101100000101001010111101010000000110000010000011010111111101111100110011000011111001001011001110101000110000101001110011110001110101010111101100000101111111011001101011111101101001011000110010001111010010000100101010101011000100101111111101001000111011000101110100110111101010000101010111101110010110001010101001011111110011100010110001110101010110110110100111101001111100011011110101010011110110010000001111111011111111011100100011101010000110000000000001011010100011011011100010011000111110011101010011011111110100011101000011100111111001100011001000111110101010101110101110101011010100010110011100010110101101000000110111001111000110111001011101110110001000111000001101111101111100111101101001100100000100110111010011011110011010111001010000011111101100111000101111011101101101000000010111110111101000010110101101100100100111000101011110000000100101110011100011100000110000011111100101100011001011100110001010100111111011101001000011001111101111000011101000010010110000111011000110010101110011010010110110001100111001101000001100000101011000000101111101110110001010010111110011101100010111111011110101101111011100110000001100011111101011011010101110100011010011111011110011010001111010011101111110110000110111001011111010000111100010100100001100000101100010001111101110001100101110000100011100010110100000111111010001100110110111100101110111101110101111001101001011001111100100010100001110100011111100001101011000000101110111011100001010000110010110111100100010100101111011000010100110110101111010101001010001010111000000110010110111000111111100111110010001111001100010000110101101011010000110000110000001010110101111111001001011001001001001111101100010001011000010000111101001011110001101001011001001011100000010100101001000110101101100110100100011010101100011111011101111011111101101000010110000101010101111001111010000000100000110110010100000010110111010011101101110010111001011100101110111010010010001110001000101010100111110011110100010010000100011001100001101011011100100101111111000110110001101110111101110110000101101011111011101001101000100111111101111001001010000000110111011100011010101111111110100111111111011001111011011101100111000100010011011111101001111101001101011010011010011001001001111010110101011100111010111111011011001010111011001110001011111001001011110000101011011110000011011001010010011010010101010001000100000111010011010011010111100000100011010011011111100100000000000100101010111111111110111110110100101001010010001010110010111111101000010110010100111110100001011111010010111001001110100010110000110010110011111101001011011010000111001111101011000110100110011001010001000101000011101010100010010110001011001001111001100100110111000100100110111010111001011111011100100011111111010011000011011000100110000110010001010110110011100110000010000011110001110001000100000001110011111100001011100001010111011111100100011110110111101010001011001000100101110010000001000011101100100010010110101000000011011000010111010110101001110011110101100001111100001111110011010110000101011101001111001101110110100000011100101001111111111100000011000111000010110011101101110011100010011100001100001000110011111101010111000001111000110001111000010101111000110111100101110101000110001111111000101001100000111010111100000100110100010000111001010000111011100001010011101001001111101100110111100011101011110110100110011011011010000000101010010011011000101011010011111111000111011101111111011110011111110001010011011001011001101100011111100000000110011001001100000101110111111001101111110110011011111111111111101010111101100010001010011101000011110001001100110101010111010110100010101011000100111011000100010011101001100111111010001101111000010110000100001001001101101100011011001010111000100001110110101110100100111011100000010010110111001101011011110100010110111111000101100001100001011100010110010011110111110001001010100011110100010011011100001011001101101010101110000001101110000100110000000100001110001101110101011001011001000010101011111101010001011110100110001000010101000011000111001110001100011011011001111010010000111100010011100110011001101001101100100100000011110000010011010001111111100100011111011001100001011000100100111111010010001100110001001100100111111010001110010111010001011110000111101110001101011011100101111011000101000101011001001111111010100000111001011011111111100011111110011101001100100100111011010000011001010100001000111001000111001110111001010100110011010000110100011111100101001011100010011010011010010111010001100111100000010010111111111000100100001110110001101001001010101100100101101110000000100100011110110000100000010111010111100011111111110100100011100010011011001011011011111111010010001011011111110011000011010011010101100010000001010110000000001001111010111010001011000000001000111001011010110110100111000100010000010010110001011111011111000010011100110010100111001111110010001010101000111101100111011010010101101101100100100010100010110101010111001011011011011010110110001101010110010000011101100010000100001011000010011111011110100110001010110100100110011010101000000010000110101111100001001011011011111010010100011010111010100000100000110101111000001000001010100100101010011001001001101011000111011101100011010011111111000100100000111010110000101100010100000010101000110111101001010111111111101011100001110000101101100010000111101110111100111010011011101100100111010100101101010111100000000110111111100110100011010111101101100100011110010101110010111110110111011100011101010101010100110110101100011111011000001110111111000100110001011100110010110011101110101101101111010111010101100101011110001111011101011111110000110001100110101101100101001100001100000010001010010001111011110010010101101010011110011101101111100011111011110101010111100110001011110101101001010000011000011000110110100110001110111001001100000011110001100111101100101111000111001110100000011001001010010110111000010110010011001110001101110101000001110011010001111011100010011000101110100001101111011111111111001100000100111110100100110100000111000110110110010110000111011111100001110101011001111010010100010111101100110001010101100100010011111011010000010010111110110100101101100110111001110000010011010111101101011010001001011001100111110001101011101010001111001010011100010011110111101010110110010101101111010011110000010000001110001110010011010111110111001001000100001111111000011000000000111110001000011110010010001110101001111001010100001011011011111010010000110111110100000101100101001111110000111011001111010100000111100100001011110101000011010101100101011011011111110110110000110011100110010100010110010111001000110001010101011100010001001111000101011100011110101110010111011001101010011011111000101011101001110101111110001110000011011000001001011110100111000001010011001100001101100001100101000110010100110001010011110001111000100001011100010011110010101111101010111101000001001100011100001001110011100010111010001011001000110010110011100100000000100100100110010110000100111110111000011010001001001100100111100011111001001100011101001111011111111100100100101011101110011001100011010111011011110100011110100010000110000100001101000100111100111010010111011111000001110000110110101111000110110100011110001100101100101000100110011011010000011110111001100100001100010110010000110101100100100010011001111010011100001011010000101110110110101101110100011001000101011010111000111000001000001110111110101101111100001011011111101111010111101000001100011101001110011100100011010001011101110110111010010001111111100101001101111111010000011001111001110110010101100101011111111110001011011110101100010110100010100100011111110010101010000010100000010000000011011111001001011111000110111110000100111100011000101100000011101011100100001111100011110000011110000001001000001100000011111000111100110010001111100111011101101110101101101100110110100001011010101101111100101110100101011100100001101111100110000010011011011001010011000001001101011010010100111001101110100001110011100100010110001010001101111011011001010101000010010001010011110110010101101110110011110101101000111110011010010001000000010100101001100110101001000001011001100011001001100100111100010100011011011100111000100000010011111101110011100100000110000110101000110011010101001010001011111010000110001010010000010100110010100000101001101111000000001001011111100100011110001101000111101000001111110110101001110000010110000000011101110111010101011111110001110110001111110101110111100011100101001000111000001001000110111010101010101101101101110110000101010010000101010001001011001110011001111011100101110101011000110010001000101000101100010011110010010100011101101110100101111000110000101111010110111011011111000111011001101101101000111100011000000101111101000001110001000000111001101011011110111110111011111001010110100000010101100011010001001110001110111111000100010010111100011011101111001001111101000111110111110100010010010110001001001011101010010001111000011101100001010000101100111001001000001010000001011111001011000111000110010100100101100010001000111100001011001011011011010011110010011011000001110011000100000010011010111111110011110010100111010101100010101101000110000010010011110001111001001111111101010010010010100011011011110000010000110110101111101111011101010001010110001011101001011000010010101111000110000100101110010100111110010010011000011111011000011010001010110100101001101010011000100011100001010000000110111001101011100010001100111010000110001000011011010100101110011000010010111111011110111011000000111011100110101110110001001110111001101001110100000100110101110101100011101100111010000111001110110010101010100011001110000110000111011000011000011101110100101001111110101101110111000001010111001100000010001001101111010000011001001001001011001110100100011000010001111011110011111010100001010110011100011010110111001001111000010110101000010110010000000000110100100001100110000111011101101000010101000100000011001011100010110100111011101101110101111100010001111000000111110110011011100011110011111010111010101000100001111010011011010011011001110001000111101100001111111000011110111010100111010101101001100111110010010000011000111011101111100000111001010011111101100011100011100001000100110011001001111000000100011110111010100111111111111111110010101100100100111001111011011011001111011011101111011100110011011001111000110000011010110011111010100101010101110011010011011011101010101011001110010000000001000000100111011010101000011100100011101001011001001100000110000101100111000100001101110000110000100111110000101110100001101100101100000101111001000001111001101101010000000111000000011010101101110101000101100100111010100010111010010010110010100010011100001011111111000010110111111010110001111001101101010001010110101110100100100001011000000110111010000011111000001101011000100101110111000100000011000011110100001100001000100010010000100100000111110111110001111001000011010001111000011110100011000010100000101110111011111001101101010010101000011111000110101111110100100110010100000110001110001000010111110001001001101000010011110100110010010111010111011011100111001101101001110111101101010101001111101111101011011011101101001111111101100001111100001011101001011101110000010101011100101100011100100001011101111011101101111101111101101110101100011101100111010001110000111111111000000001001100101001011010010001011010100110000001011011010001001010100000100110011011011100010011100000001111101101110010001010110101100001101010101011100000001100011111101110001010000011001010001100001010001011000100100010110000000001010001110000010111110111101110100010110001101001100011001101111101011111110001111100100111001111111010010011111110100100000100101011001010011100110010010001110110101100111101110011100101100110110111001001011111101111100101001110101110110101010001110111111010011010011100110100111101110010111011011001000110111110000110111101001111011101100110000111010111011100000000010101110000100010100001101001011010011010100011000110010000000010111001001101100101100111101000111011010110100101101101000010101011000100011011100010100101101101100010001101011101011100111001011010010001100101011100111111000101000111010110110110000101000000001101100000110111011101011111011101010101101011100001010111100000100011000010101101100001011111011110100011110001111110110001000111000100001001010000001111101111011100101110101001100100100110111100110101000000100100101000101010001110000010111110110010011111011110000011100111110011100100111101000110010110000100110110111101110100001110111001111010000110100010101011001100011001100100010101110111100000001100111000111001000011100100101010101101110011000100100111101011101100110010001111100001110100110001111010001000101110011001100010001111001111110110100100011111101101010100000001000001110100101010101001111111100100000101111010000101110010010001000011010101110001000001111100100101111011111010110110100010111110110011011001010010000001010100110010101100010000001100010111101100110001010001101111111000111101010011101000011000001001110110110100001111000110100111011010000101010101010100101110111011110111110111100110010010001000010001001111110101001001010110110000011000100101010100101000011011111011011011100011111110001111001001011110110000111001011100100110011110000110000110111001011011000010101011011001000011010011110111010101100010001101001000001111010011011111100111100111100110101111111110000110001110000100111011000010111001010101100100110000110011010011100110110111000100111101101111101001111001001101100000000110000000110001101000100000011110010010101110110100010001011100100011101011010000001111101001001000101001011000111011100011101001010010000111010010111111100111111111001010001110011010110001101110010110111010110001101111100000111100010101100000111001000011110100001000111100011111110000101110010110111011010000001010000001010111011100011011011000000010100110001101110000101110011001010011000111111111101111001001101110111111110001001110001111100111100011010101110011101100000010111100111010011000011100010111101110100111011000110011001010011000100011100000010110110010011000000111001011010001000101101100000111101110100010100010010100110100001001101010111011001001100101111010100010000111101001100110110010111001010100100011100111001011000010100111100010110100010111000010101100110001100111111111100011111111000110110000110001100000111000011001010100010110001110001011011110111001010001001001010010010011101000010111110011101110110000110001001101111001001100100111111011111010100001101101000011100110101111000011011010000000111000011011001010101101101000001011011101101010101000011101011111001000100100001010010000101010111010000101000110001110100101110011001100010110000110100000110101010110100010011100000010001001000101100101111111111001011011101010110101111100110000111000111000111111100010011001000010100100101001110010101001101110010001110111000000011011101110011110100011100100010001110011100100000010001110000010111010110101000111111001110111111111000100001011000000011010111100100111011001111000001000101101000111001110110111000010010111000000100101010001110011101101011010010110100000100100111000001011110011010000001111011010101110001010110110100110001010001001000001001110100111010100101100111110101100011111100000110000101010100010000000010001000010011001100101000101000111011101100100000000100101101011110001111010000111001100010101011101110001011111110110001010111011011010110100100111000101110111010100111100111010110011001000110011100100010001010001111011001000100000110101100010111010110111110011011010000110100101111000010000010010010100100010000011000001111111010000010111101101111111111000001011010000100101001000010100011001000011111110101111110011011010110101011100001110101101100001010100100100100010100010111001011001001000100001000101111100110000101100011101111110111001110001100100101001001110101011001011001001110101011011010001011110001010001010001101111000101011011011010001100011010101010100001100001010010001101001010001101111101110001110000001110000000100100000101001011010100100100001010100010000001000000011011111110001110001011011100110110010011111111001001001011011011110010010000110111110111011101110000010100010110111110010111001110000010010001111100011001000101001111011100001000101100001011110010000111001111000000111000101101111000110010011010011011001001000001010000101100001100000010011100010100000010111101101011110000101111111011001001111101010000010110011100110101110001001110100000100100101000010011100100011010111110011010000011100100111010011011011010100010111110011001010011100101000001100111001101111010111101001100001010010010110101000011101000110100111010001011011111000110000011110101011010010101000100101011101011111010000110110010100000011111001101111100111010111010001001010111101011001101101100110001011100100110001110110000011010011000010110010100001001101101000110001010110100100100101011000110111011100110100000111110000001010001001010100100101001001010010100111010111110100100001000010010111001000101100010110100011110000100001011001011101110111111101000100101001001101000101000010000110010110010010110011000011111011011000001101000111100000100001010111101011000100010000001110100111011100001010001110010001100101111000110001000000110101100110001010010111000000110011110011101001011011100011111001111110110001111101100111011010100000110111001101000111010110010111011100000001010110001010110111100111101010001110110100010000000010101101101011011100011100000111101000010001011110100111001011101111101110001111111011001110000010110101001101011110110001101101110101111000100011100101010100111110001111000000001111101001100011001001111101111011001101000110111010001111000100011100100000010001011001100000000100010111010101010101010100111101100001010110000001101111101101100110001010011000110001100110111110110101101001001100111100100100110010110101001100001101101110110100110110001110000010111001111111100011101001100101001101111110011011010000101110110100110111111110001100100011011111010111100100101101110101010111000111101000101000110000100010100101101101001011111100010000010101101110101000100011101101011110010001110001010010100000101000011101111011100100110000110110100001001001100100010101010010101001100010110011011100110111101110100011111010111111011111110101100000011010010001100000110100111110010100101000011101000010100110010110001110000000000101110011110010001010011100001101011100100000110000100101101000011110101010110101110110110001111011100101100100101100010000101101010100110111010000000111100100110000110111110001110101110100011110010011111100010001101010010001100110101101101001110110000011000000011001010110000000110010011101110001011010100010100111100010001010010011101010111101001101011111011001010001010011011011111010001110011011111010110001001001011000101000010000001001000101001111110100000011100110000001111010011101000101111001001111100101100100010011011001011100010011101111010111111110001111011000111111011111011111010100001001011011101110001011010110111001010111101110001111000110101000110101000110011101110101110111010110101101000010000110101110001010111010000001110110101100111001011100110110011001110010001011001010001000110011111011010000000011101010101011111011001011101101010010110100110111010100000100111011000100011101000011100100100110111110001010111010111110011000000010110100000101111110010101111100011000111001001011001010000101101010111001000000100100100010000111110111011101100111010001011011111111101000001111011010111011100101001100100111011101101000001001001010011010010100010011100000110000001001001101001110000101000010100000010111111100111000001011000111001110101101111000010011111011010100011101010001100101010101101011101110001110010101011001001111101100101111011101110000000111000111101000111011110010111000101011100100101000111000011101000001100001111001111111001010001010011011111111001000110010101011000101111000011001101100011111101000110001011001000010000110011010000100010101101101001011001110111010101011001111110011100110111110001100011110001111001011010010101111001100111101010011100000110010000100110101011111111011110110010111011101111100011111110000110010101001001100010100010111000001010010011010011010111110010001010101011011110011110000001010110101101010001001000110111110111110110001100000000011110010010010011011110101011001011010101011000010011010111100000000111001000100110011101000111101001001001101101110111101100100011011001001101110011001101000011100001011010001111101010100000110001110101101101100011011011110000100010000110110100111100111011010001110100000101110011110110100101100010110010101101010111101111000101100110011111010001110000111010110001010110111110011010001101111110000100011001010101010101101011111001001000000100011001110101000101110011001000100100011101110100000110111111101110000010010101011110001011111101111110101110101100110110101010100101001010101011011001010000000110110000101110100010011011011010111100000001101011010111100110010101100000001111100100100110001111011000001000110010100011111010010000110000110011101000110110111110011011001101001001101110011101101010110000111010000001110010110101011000100001011000110110000000111100110111100001000000110111001011100010100001111011110100001010010010000010110001011110101010110011010100100001110101001111010100100110010101111010000110100100101111011111100011000101101010101110001010011100101110011111000100110101101101101001110111110100100100110010010000010001100000011010010110101010001100100000010001001110010111010110101010101110011110101011101010010111110000111001010100010101001001011000111011010100100100011110111011011101111110001110110000010011011010110111100100010111100101010111000001100110110101101101100011001011010010110000110101010111000101001000010011101011110111000011001010110000001001111110100110011110010011101111111111010111011010111111101010010000011000000111011010100010101010110101110110110001001001111010010010001000001100111101010000011001101111011111011101110000100000011011110001001101010111111000001100101101000000111100100001000010100011101011111000110010001111010001011001001111000011011111100011011111001100001011011100001100111111011111001010101011111011001010011111000111001001100000001101010111110000101011010011111100110011111101011111001100101101101101010111000011110011111010010100011111001110111011010100010111011001111111010100011101001000011001010111111110110111000001101101100111111111111111011110100000110011111001010110011110111010100011110111111011110010010101100000000100011100100000001000101000100110011100100001000011001111010101110101101001000110111001101011000100110101000111111110101001100111000011000100101110101100010100000001111111010011001010010001001010101011101110000010011010000000100110011000010000000110111000101001010101110100110011100000101111111001000010111110111010000110110110001100111001010110000010111001000011101111011010010111100011110111011111101001000111000001101010001111110100110000011011001001011100101101101110100100011010011111101111001001010101101000011110001011111001100111010101100010011011001011110110000110011010111110111011111101111101000010001000011101001100110100011101000111110101111110111111110000110000110111010101010011011011100110000110111011000010000110000111001011111001001011001100101011111000001000000011000110100010001011011100010110101011000101110111101101010101100111101000000110011110011110110110110110100000100010010000011000011110000010000001101000100100000011010001110010001000100010010011000110000011111100101010010001111111000111101000100100111001011011011000011001000011101100011110100011111110111011100000001000100111000111001110000011100100011110001010010101100110000100100010000000110110010110000100001101111011011010001010001100001011111110111010111011100100000011101111111101110111101001100001101011010100101010010001000101001111010011101100011110111000111010000010100010111001000101101100010111101111010110111110111111001100100011011000111100011101011001101010110111100010100000001001000110100100110100010100000001001010111110111000001101100101111011000100100011010111000010000100010001011110011110010111001000111001101100101111001000101110100011010000011000000110110111100011101101100010000101000111101100010001110000110001010100111000100011011101011100111001101110001110100111001100001011001011000111111111111110111110101101110100110000101100101101111000011100111011101101000101111110000100101011001111101101001110001010001110011001100000001111101100110001111111101100010101110011011001110011010110111001000001110111011001001101110010001000111001001011110110011101100000110010000111111101101011010111011100010101001011110101111011111100110111101011111100101100100000110100000100101101000000111110100011110011101011000011010110110111101101000000111111100011011011010100101100001000010001101101101111011001111001110111010111101100100100011001010110110111111011100010101001000100011001101000001110001101011011010110111000111001100100111001110010101111000100101101000011011001000010101101110011100001000111000110111011101011010001100111000110110101111110101000010011110011000110001000001010100001100100001001110001101111000001111011111001100100100001010100110111000110111110100011110011001011001100111010100010100001001011111000010001010011011000011111001001110111011000011011010100110011110111011110111111111010111011010010111110100110111010000010011100110000111101010011111110010100011101101111001100111100011000001010111011110110101001111010011100011001101100000110111110100110110101110100000011101011101011001111111010100101100100010000111110000111011111101101011010111000000111100001010000001010101111111011100111001001010000000001011000011010110011001011101000011011111010110100001111100101001101101101110110110001110001000111010001000100001010000101110010111001001111001000111000110010001010010001010";

	TYPE registers IS ARRAY (0 TO N_EVENTS - 1, 0 TO 3) OF INTEGER;
	SIGNAL registers_check : registers := (
		(0,187,0,0),(84,187,0,0),(0,0,0,199),(36,0,0,199),(36,0,0,106),(0,197,0,0),(0,254,0,0),(0,254,205,0),(0,254,205,10),(0,154,205,10),(0,154,116,10),(0,154,116,242),(0,154,233,242),(82,154,233,242),(82,154,233,197),(82,154,233,213),(82,236,233,213),(136,236,233,213),(136,7,233,213),(149,7,233,213),(149,7,89,213),(149,7,89,109),(149,7,167,109),(149,7,72,109),(149,7,11,109),(149,124,11,109),(149,124,11,183),(149,124,202,183),(149,124,227,183),(149,124,100,183),(149,124,100,78),(149,252,100,78),(149,239,100,78),(149,239,100,65),(149,27,100,65),(149,156,100,65),(166,156,100,65),(166,156,85,65),(132,156,85,65),(0,0,0,95),(0,27,0,95),(215,27,0,95),(215,27,64,95),(215,185,64,95),(215,69,64,95),(10,69,64,95),(189,69,64,95),(189,69,64,109),(28,69,64,109),(28,237,64,109),(28,237,60,109),(28,81,60,109),(28,81,38,109),(233,81,38,109),(233,81,127,109),(233,81,127,235),(183,81,127,235),(183,214,127,235),(183,155,127,235),(183,155,14,235),(183,155,14,133),(237,155,14,133),(20,155,14,133),(247,155,14,133),(247,138,14,133),(160,0,0,0),(197,0,0,0),(197,244,0,0),(197,244,35,0),(154,244,35,0),(154,80,35,0),(154,80,35,65),(189,80,35,65),(150,80,35,65),(150,80,206,65),(150,80,206,167),(150,177,206,167),(150,177,194,167),(150,177,188,167),(150,177,59,167),(150,177,53,167),(219,177,53,167),(0,234,0,0),(0,234,0,204),(0,239,0,204),(0,239,0,97),(120,239,0,97),(188,239,0,97),(188,190,0,97),(0,0,185,0),(0,123,0,0),(0,86,0,0),(0,228,0,0),(0,117,0,0),(192,117,0,0),(192,117,148,0),(0,85,0,0),(0,0,0,23),(79,0,0,23),(166,0,0,23),(166,190,0,23),(166,190,203,23),(166,190,203,145),(111,190,203,145),(81,190,203,145),(81,190,203,16),(183,190,203,16),(183,190,61,16),(183,190,61,228),(183,190,61,99),(29,190,61,99),(29,190,152,99),(29,215,152,99),(29,215,41,99),(29,215,237,99),(29,215,237,214),(29,215,203,214),(29,130,203,214),(29,130,165,214),(29,130,194,214),(29,130,166,214),(29,221,166,214),(29,41,166,214),(233,41,166,214),(233,41,166,36),(0,254,0,0),(0,254,0,85),(0,254,0,72),(0,42,0,72),(0,57,0,72),(0,57,221,72),(0,32,221,72),(0,32,81,72),(0,38,81,72),(7,38,81,72),(7,38,81,27),(7,38,57,27),(7,52,57,27),(148,52,57,27),(148,52,115,27),(148,60,115,27),(162,60,115,27),(162,60,74,27),(162,60,61,27),(162,60,17,27),(16,60,17,27),(16,131,17,27),(16,131,191,27),(34,131,191,27),(34,131,191,165),(241,131,191,165),(13,0,0,0),(13,0,0,238),(160,0,0,238),(160,0,0,55),(24,0,0,55),(24,0,0,171),(24,0,0,202),(37,0,0,202),(37,0,0,135),(37,76,0,135),(139,76,0,135),(139,71,0,135),(0,0,66,0),(156,0,66,0),(0,0,156,0),(0,0,156,0),(0,64,156,0),(186,64,156,0),(186,64,156,173),(186,64,156,151),(186,50,156,151),(186,50,197,151),(186,50,103,151),(186,208,103,151),(186,146,103,151),(186,146,103,155),(186,146,103,105),(84,146,103,105),(197,146,103,105),(197,250,103,105),(197,250,103,40),(197,250,103,129),(197,250,144,129),(197,250,144,17),(197,250,7,17),(197,250,7,170),(197,180,7,170),(197,180,7,68),(197,180,154,68),(0,122,0,0),(151,122,0,0),(39,122,0,0),(39,0,0,0),(0,66,0,0),(0,66,0,27),(0,66,0,148),(0,167,0,148),(0,167,0,63),(0,0,164,0),(0,0,82,0),(0,0,72,0),(0,0,152,0),(0,0,152,185),(0,0,45,185),(0,204,45,185),(0,204,45,245),(0,0,0,4),(0,0,65,4),(0,0,211,4),(0,116,211,4),(0,116,242,4),(223,116,242,4),(223,70,242,4),(79,70,242,4),(79,70,85,4),(79,70,23,4),(79,52,23,4),(79,191,23,4),(170,191,23,4),(170,191,178,4),(170,111,178,4),(170,111,178,250),(40,111,178,250),(0,0,176,0),(0,0,176,91),(0,51,176,91),(0,51,212,91),(0,137,212,91),(158,137,212,91),(92,137,212,91),(92,137,217,91),(76,137,217,91),(76,137,217,185),(76,11,217,185),(76,11,217,175),(76,11,217,17),(76,204,217,17),(76,204,217,103),(0,0,0,228),(0,0,48,228),(215,0,48,228),(215,0,59,228),(215,0,59,19),(215,0,0,19),(215,0,0,4),(215,0,0,105),(199,0,0,105),(97,0,0,105),(97,0,74,105),(97,0,65,105),(97,0,65,207),(97,155,65,207),(97,155,90,207),(97,83,90,207),(97,83,90,124),(97,113,90,124),(97,217,90,124),(97,106,90,124),(215,106,90,124),(21,0,0,0),(134,0,0,0),(134,185,0,0),(57,185,0,0),(57,185,243,0),(0,0,87,0),(0,0,75,0),(0,0,227,0),(0,0,38,0),(68,0,38,0),(50,0,38,0),(0,7,0,0),(107,7,0,0),(137,0,0,0),(137,0,0,245),(137,137,0,245),(137,155,0,245),(137,155,248,245),(17,155,248,245),(81,155,248,245),(22,155,248,245),(22,150,248,245),(22,150,178,245),(94,150,178,245),(94,150,178,233),(94,150,1,233),(94,150,101,233),(94,150,101,84),(0,0,0,253),(0,0,98,253),(0,0,98,207),(0,206,98,207),(0,206,34,207),(0,206,34,182),(0,206,114,182),(0,206,240,182),(0,88,240,182),(0,214,240,182),(0,172,240,182),(196,172,240,182),(196,172,151,182),(196,172,7,182),(196,172,202,182),(196,172,202,1),(172,172,202,1),(172,172,244,1),(172,172,244,27),(172,34,244,27),(0,0,64,0),(0,0,37,0),(124,0,37,0),(124,0,37,213),(124,0,224,213),(0,0,0,245),(0,0,0,205),(0,56,0,205),(0,56,80,205),(0,56,80,255),(0,56,146,255),(0,56,146,96),(0,107,146,96),(0,107,199,96),(0,107,88,96),(21,107,88,96),(21,39,88,96),(21,39,206,96),(21,39,206,199),(21,39,144,199),(21,39,158,199),(21,46,158,199),(0,207,0,0),(0,207,153,0),(0,109,153,0),(0,133,0,0),(0,133,148,0),(0,133,148,127),(0,133,148,67),(0,98,148,67),(0,240,148,67),(0,58,0,0),(0,97,0,0),(9,97,0,0),(9,2,0,0),(9,2,67,0),(9,2,127,0),(9,2,127,229),(9,2,127,20),(0,0,10,0),(0,0,116,0),(0,105,116,0),(0,166,116,0),(0,5,116,0),(252,5,116,0),(220,5,116,0),(172,5,116,0),(172,5,116,179),(172,5,116,65),(172,5,147,65),(172,5,147,68),(172,5,21,68),(172,5,21,203),(194,5,21,203),(76,5,21,203),(76,11,21,203),(76,121,21,203),(0,0,85,0),(0,0,85,33),(211,0,85,33),(211,0,193,33),(211,223,193,33),(211,91,193,33),(211,91,193,210),(211,91,19,210),(119,91,19,210),(104,91,19,210),(28,0,0,0),(28,0,0,178),(28,0,23,178),(28,0,23,218),(28,90,23,218),(28,90,23,182),(28,229,23,182),(28,229,23,90),(104,229,23,90),(104,120,23,90),(251,120,23,90),(0,0,0,144),(0,132,0,144),(170,132,0,144),(170,226,0,144),(170,226,0,212),(0,0,0,247),(0,0,0,61),(0,236,0,61),(0,156,0,61),(27,156,0,61),(86,156,0,61),(86,174,0,61),(86,86,0,61),(55,86,0,61),(55,115,0,61),(19,0,0,0),(19,0,111,0),(19,0,200,0),(19,0,236,0),(19,0,226,0),(19,0,37,0),(19,0,37,185),(19,0,173,185),(19,0,194,185),(19,0,104,185),(101,0,104,185),(101,20,104,185),(101,20,104,35),(101,20,104,110),(101,196,104,110),(101,174,104,110),(101,174,104,88),(101,221,104,88),(101,221,104,33),(101,221,104,112),(101,254,104,112),(101,254,104,226),(101,254,104,226),(101,130,104,226),(101,181,104,226),(101,181,104,177),(101,181,104,157),(101,181,104,12),(0,0,0,194),(0,0,14,194),(0,168,14,194),(0,0,0,194),(205,0,0,194),(205,229,0,194),(205,229,215,194),(205,240,215,194),(205,240,215,132),(116,240,215,132),(116,240,215,215),(116,142,215,215),(116,215,215,215),(116,161,215,215),(135,161,215,215),(141,161,215,215),(0,0,216,0),(0,100,216,0),(0,0,0,193),(0,0,202,193),(0,0,36,193),(0,0,58,193),(0,166,58,193),(0,166,58,93),(0,166,58,131),(118,166,58,131),(118,203,58,131),(118,154,58,131),(118,118,58,131),(118,118,228,131),(118,118,228,235),(118,118,249,235),(118,118,249,126),(118,7,249,126),(0,0,0,73),(174,0,0,73),(174,0,55,73),(20,0,0,0),(70,0,0,0),(70,151,0,0),(27,151,0,0),(27,151,14,0),(0,0,140,0),(0,0,171,0),(0,0,171,244),(0,53,171,244),(214,0,0,0),(246,0,0,0),(246,0,0,54),(246,0,13,54),(246,169,13,54),(143,169,13,54),(54,169,13,54),(54,169,13,44),(54,169,13,69),(54,169,1,69),(54,90,1,69),(54,90,158,69),(54,90,158,116),(54,90,88,116),(54,222,88,116),(54,222,172,116),(70,222,172,116),(70,222,196,116),(70,131,196,116),(70,131,196,189),(70,131,65,189),(70,44,65,189),(185,44,65,189),(185,44,65,241),(185,44,65,120),(185,44,136,120),(185,44,123,120),(185,99,123,120),(185,99,123,42),(185,99,10,42),(185,99,10,204),(185,219,10,204),(129,219,10,204),(129,37,10,204),(129,175,10,204),(241,175,10,204),(19,175,10,204),(169,0,0,0),(171,0,0,0),(171,73,0,0),(171,73,0,164),(58,73,0,164),(58,73,80,164),(58,73,80,84),(58,61,80,84),(58,152,80,84),(58,152,80,13),(58,143,80,13),(99,143,80,13),(158,143,80,13),(158,143,80,194),(158,143,80,32),(158,86,80,32),(158,86,120,32),(158,86,120,191),(158,86,128,191),(158,187,128,191),(158,187,187,191),(158,187,33,191),(247,187,33,191),(75,187,33,191),(75,187,33,159),(114,187,33,159),(144,187,33,159),(0,96,0,0),(0,196,0,0),(0,196,0,99),(0,196,183,99),(140,196,183,99),(244,196,183,99),(244,196,216,99),(244,47,216,99),(70,0,0,0),(70,0,0,163),(70,0,163,163),(70,0,163,84),(66,0,163,84),(66,202,163,84),(66,202,64,84),(66,202,64,125),(66,202,131,125),(210,202,131,125),(210,51,131,125),(210,150,131,125),(225,150,131,125),(225,174,131,125),(0,0,0,10),(195,0,0,10),(0,0,0,94),(255,0,0,94),(185,0,0,94),(185,0,0,212),(208,0,0,212),(208,251,0,212),(134,0,0,0),(24,0,0,0),(24,0,51,0),(21,0,51,0),(97,0,51,0),(45,0,51,0),(54,0,51,0),(15,0,51,0),(132,0,51,0),(132,121,51,0),(132,114,51,0),(86,114,51,0),(86,114,51,19),(30,114,51,19),(30,114,51,85),(30,114,227,85),(156,114,227,85),(156,114,227,236),(156,114,201,236),(156,114,201,154),(46,114,201,154),(159,114,201,154),(198,114,201,154),(198,114,201,184),(118,114,201,184),(118,114,116,184),(118,114,252,184),(118,114,252,183),(0,0,164,0),(0,97,0,0),(0,97,0,152),(0,6,0,152),(0,6,0,23),(0,6,213,23),(0,6,213,9),(0,1,213,9),(0,1,213,198),(0,1,213,102),(0,1,90,102),(0,1,57,102),(58,1,57,102),(58,61,57,102),(150,61,57,102),(150,61,57,36),(199,61,57,36),(199,61,57,99),(142,61,57,99),(31,61,57,99),(31,61,57,88),(31,61,167,88),(0,40,0,0),(0,40,155,0),(0,40,206,0),(0,176,206,0),(0,123,206,0),(0,123,206,122),(48,123,206,122),(48,123,189,122),(48,123,189,99),(0,0,0,44),(29,0,0,44),(0,120,0,0),(0,26,0,0),(0,196,0,0),(119,196,0,0),(119,196,69,0),(178,196,69,0),(178,196,69,11),(0,0,0,4),(0,0,0,109),(0,0,105,109),(0,193,0,0),(0,193,0,113),(0,193,0,45),(0,0,0,49),(0,0,0,116),(80,0,0,116),(80,0,0,243),(152,0,0,0),(152,0,0,31),(152,126,0,31),(2,126,0,31),(0,0,105,0),(0,1,105,0),(0,1,105,204),(0,1,105,70),(0,1,150,70),(0,1,150,56),(0,1,150,194),(0,1,150,70),(0,1,150,130),(167,1,150,130),(167,96,150,130),(167,96,169,130),(203,96,169,130),(203,96,169,167),(203,150,169,167),(203,150,222,167),(223,150,222,167),(223,150,186,167),(83,150,186,167),(83,66,186,167),(253,66,186,167),(253,185,186,167),(253,185,2,167),(253,145,2,167),(139,0,0,0),(139,139,0,0),(139,60,0,0),(139,60,0,106),(139,95,0,106),(139,125,0,106),(195,125,0,106),(195,80,0,106),(195,80,0,56),(195,126,0,56),(195,126,0,91),(175,126,0,91),(2,126,0,91),(2,126,0,12),(2,126,0,70),(73,126,0,70),(73,126,0,27),(157,126,0,27),(157,126,83,27),(123,0,0,0),(123,203,0,0),(123,203,0,218),(0,0,39,0),(0,96,39,0),(0,96,0,0),(0,96,198,0),(0,96,139,0),(121,96,139,0),(121,96,139,40),(121,96,139,181),(121,96,139,14),(121,96,183,14),(121,96,183,49),(121,96,232,49),(121,96,232,164),(193,96,232,164),(193,96,168,164),(230,96,168,164),(230,114,168,164),(230,114,222,164),(230,109,222,164),(230,107,222,164),(195,107,222,164),(195,107,222,60),(0,0,165,0),(141,0,165,0),(141,0,230,0),(141,0,166,0),(141,0,21,0),(141,252,21,0),(141,248,21,0),(141,248,181,0),(141,248,72,0),(225,248,72,0),(225,64,72,0),(225,64,72,75),(225,64,19,75),(0,0,0,84),(146,0,0,84),(146,0,0,51),(88,0,0,51),(88,0,98,51),(88,0,5,51),(177,0,5,51),(177,0,193,51),(57,0,193,51),(57,0,89,51),(57,83,89,51),(57,83,15,51),(0,0,0,121),(0,82,0,121),(0,82,0,177),(0,85,0,0),(188,85,0,0),(188,85,224,0),(188,85,53,0),(70,85,53,0),(70,85,53,158),(70,146,53,158),(124,146,53,158),(124,146,53,243),(213,146,53,243),(213,13,53,243),(213,13,178,243),(213,13,178,37),(0,0,2,0),(238,0,2,0),(238,0,2,99),(238,0,2,158),(238,0,2,145),(238,0,2,49),(238,0,2,206),(238,0,60,206),(207,0,60,206),(207,113,60,206),(207,113,104,206),(123,113,104,206),(123,113,104,169),(123,113,142,169),(123,238,142,169),(123,129,142,169),(0,0,92,0),(0,0,113,0),(0,89,113,0),(111,89,113,0),(177,89,113,0),(177,212,113,0),(102,0,0,0),(102,0,0,7),(102,0,118,7),(0,0,57,0),(0,0,224,0),(229,0,224,0),(229,199,224,0),(229,199,255,0),(229,199,25,0),(229,199,25,19),(229,177,25,19),(229,134,25,19),(0,16,0,0),(0,11,0,0),(0,11,0,248),(0,93,0,248),(0,93,129,248),(0,125,129,248),(0,29,129,248),(100,29,129,248),(100,29,228,248),(0,205,0,0),(0,205,0,103),(0,205,235,103),(0,205,126,103),(0,205,94,103),(0,205,94,218),(0,131,0,0),(0,131,0,59),(0,141,0,59),(0,239,0,59),(145,239,0,59),(145,239,0,222),(0,172,0,0),(0,199,0,0),(0,163,0,0),(0,253,0,0),(0,253,212,0),(0,250,212,0),(0,250,37,0),(0,250,37,0),(0,250,220,0),(41,250,220,0),(41,250,3,0),(41,250,247,0),(41,250,21,0),(0,0,113,0),(0,0,197,0),(0,0,216,0),(0,0,216,38),(0,0,41,38),(0,46,41,38),(0,46,41,189),(0,222,41,189),(0,247,41,189),(0,247,41,19),(0,247,41,249),(0,247,41,179),(0,247,143,179),(204,247,143,179),(204,13,143,179),(204,13,91,179),(243,13,91,179),(0,0,139,0),(0,8,139,0),(0,225,139,0),(246,225,139,0),(246,225,139,77),(0,0,193,0),(0,0,193,201),(0,0,167,201),(0,117,0,0),(0,117,0,141),(0,67,0,141),(162,67,0,141),(0,0,73,0),(141,0,73,0),(141,0,73,0),(141,0,179,0),(141,0,140,0),(210,0,140,0),(0,0,0,46),(0,206,0,46),(0,186,0,46),(0,186,10,46),(0,186,58,46),(0,129,58,46),(0,129,58,46),(0,129,2,46),(51,129,2,46),(0,105,0,0),(212,0,0,0),(251,0,0,0),(251,0,69,0),(251,206,69,0),(251,206,69,60),(251,206,69,120),(251,64,69,120),(251,64,69,131),(251,64,235,131),(31,64,235,131),(31,197,235,131),(31,209,235,131),(0,0,52,0),(0,0,52,135),(0,47,52,135),(0,47,215,135),(44,47,215,135),(44,47,173,135),(0,0,191,0),(0,0,104,0),(0,12,104,0),(0,90,0,0),(0,90,0,28),(0,0,0,39),(0,219,0,39),(0,219,181,39),(0,96,181,39),(123,96,181,39),(212,96,181,39),(212,96,181,79),(212,33,181,79),(212,208,181,79),(212,165,181,79),(212,165,59,79),(0,0,0,79),(0,0,128,79),(0,0,0,30),(0,0,0,172),(168,0,0,172),(168,0,0,237),(168,0,92,237),(168,0,92,138),(168,104,92,138),(168,133,92,138),(168,133,128,138),(168,133,128,225),(147,133,128,225),(147,133,128,141),(31,133,128,141),(31,133,128,195),(31,133,128,138),(13,133,128,138),(13,133,128,15),(13,133,128,105),(13,37,128,105),(13,37,157,105),(55,37,157,105),(55,54,157,105),(0,118,0,0),(0,118,0,146),(0,118,117,146),(0,118,117,85),(0,118,117,53),(0,118,161,53),(0,118,161,153),(73,118,161,153),(73,176,161,153),(73,176,161,49),(73,203,161,49),(153,203,161,49),(9,203,161,49),(160,203,161,49),(0,0,159,0),(252,0,159,0),(252,0,39,0),(252,0,39,18),(107,0,39,18),(0,0,0,142),(99,0,0,142),(0,74,0,0),(0,74,206,0),(0,74,206,216),(0,74,174,216),(0,213,174,216),(0,213,174,31),(0,151,174,31),(0,151,199,31),(0,151,199,12),(133,151,199,12),(133,219,199,12),(133,219,199,248),(133,219,199,149),(133,219,199,1),(220,219,199,1),(220,219,199,39),(220,219,142,39),(220,219,142,50),(220,219,142,236),(220,219,244,236),(22,219,244,236),(22,21,244,236),(25,21,244,236),(179,21,244,236),(179,21,176,236),(0,252,0,0),(0,251,0,0),(0,8,0,0),(180,0,0,0),(180,105,0,0),(187,105,0,0),(0,0,0,38),(0,0,118,38),(0,0,118,132),(0,0,217,132),(0,142,217,132),(0,142,133,132),(0,142,133,44),(168,142,133,44),(37,142,133,44),(37,142,133,182),(37,116,133,182),(37,116,133,249),(37,116,133,26),(37,32,133,26),(37,32,133,165),(37,221,133,165),(37,93,133,165)
	);

	SIGNAL do_reset : std_logic_vector(0 TO N_EVENTS - 1) := "1010010000000000000000000000000000000001000000000000000000000000010000000000000000100000011000001100000000000000000000000000010000000000000000000000000100000000000101000000000000000000000000100010000100000001000000000000000010000000000000010000000000000000000010000100000101000000000000001000000000000000000010000100000000000000001001000001000000010000000000000000010000000001000000000010000100000000010000000000000000000000000001001000000000000101000000000000000100100001000100000000000000000000000000000000000011000000000000000000000000010000000100000000000001010000010000000000000000000000000001100000000000000000000100000000101000000100100100010001000000000000000000000001000000000000000000100100000000000000000000010000000000001000000000001001000000000000100000000000000010000010010000000011000000010000010000010000000000001000000000000000010000100100010000010000000011000000000001000001001010000000000101000000000000000000000100000000000001000010100000000000000000000000010010010000000000000000";

	TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL RAM : ram_type := (
		75 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		96 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		135 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		151 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		190 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		284 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		309 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		402 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		469 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		477 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		664 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		676 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		703 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		810 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		833 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		853 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		906 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		1005 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		1176 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		1243 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		1358 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		1372 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		1424 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		1566 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		1579 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		1717 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		1779 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		2003 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		2004 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		2008 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		2159 => STD_LOGIC_VECTOR(to_unsigned(18,8)),
		2176 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		2349 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		2354 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		2402 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		2406 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		2550 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		2580 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		2608 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		2637 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		2694 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		2740 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		2824 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		2833 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		2846 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		2856 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		2871 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		2915 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		3004 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		3026 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		3356 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		3493 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		3639 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		3669 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		3732 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		3789 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		3822 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		3830 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		3852 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		3941 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		4042 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		4069 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		4090 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		4106 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		4244 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		4267 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		4293 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		4403 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		4414 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		4469 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		4516 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		4521 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		4767 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		4806 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		4900 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		4928 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		4952 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		4986 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		4995 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		5051 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		5126 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		5231 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		5339 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		5351 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		5425 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		5438 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		5444 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		5447 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		5543 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		5591 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		5600 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		5611 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		5639 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		5671 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		5684 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		5695 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		5806 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		5839 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		5872 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		5896 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		6031 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		6117 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		6127 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		6134 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		6172 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		6388 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		6481 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		6727 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		6764 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		6806 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		6896 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		6933 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		6971 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		6975 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		7023 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		7147 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		7268 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		7310 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		7369 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		7376 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		7452 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		7590 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		7803 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		7806 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		7931 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		8085 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		8246 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		8293 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		8318 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		8452 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		8523 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		8545 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		8579 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		8679 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		8773 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		8788 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		8843 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		8898 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		8925 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		8953 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		9123 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		9125 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		9134 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		9173 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		9209 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		9283 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		9297 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		9326 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		9393 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		9474 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		9532 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		9614 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		9699 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		9729 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		9815 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		9835 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		9903 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		9930 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		9940 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		9996 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		10000 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		10071 => STD_LOGIC_VECTOR(to_unsigned(3,8)),
		10158 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		10351 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		10513 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		10611 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		10644 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		10649 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		10679 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		10776 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		10789 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		10827 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		10865 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		11121 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		11345 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		11374 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		11379 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		11456 => STD_LOGIC_VECTOR(to_unsigned(137,8)),
		11458 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		11482 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		11490 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		11555 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		11675 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		11693 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		11815 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		11908 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		11967 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		11989 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		12130 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		12192 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		12219 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		12367 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		12385 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		12504 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		12625 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		12644 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		12659 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		12871 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		12946 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		12961 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		12973 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		12977 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		13062 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		13089 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		13192 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		13208 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		13248 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		13380 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		13383 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		13384 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		13468 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		13484 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		13488 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		13550 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		13559 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		13578 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		13579 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		13627 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		13711 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		13750 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		13910 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		13925 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		13986 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		14104 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		14108 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		14113 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		14127 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		14172 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		14201 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		14292 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		14351 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		14548 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		14615 => STD_LOGIC_VECTOR(to_unsigned(149,8)),
		14618 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		14793 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		14949 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		15126 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		15386 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		15484 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		15508 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		15610 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		15638 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		15647 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		15944 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		16049 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		16200 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		16253 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		16262 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		16269 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		16281 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		16328 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		16351 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		16449 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		16538 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		16552 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		16679 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		16694 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		16887 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		16956 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		16986 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		17023 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		17042 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		17098 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		17119 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		17141 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		17170 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		17249 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		17348 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		17391 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		17432 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		17491 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		17538 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		17539 => STD_LOGIC_VECTOR(to_unsigned(95,8)),
		17650 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		17683 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		17705 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		17780 => STD_LOGIC_VECTOR(to_unsigned(16,8)),
		17910 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		17938 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		17985 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		18001 => STD_LOGIC_VECTOR(to_unsigned(31,8)),
		18035 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		18340 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		18374 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		18411 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		18494 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		18555 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		18599 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		18941 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		18984 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		18986 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		19004 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		19059 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		19065 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		19097 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		19258 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		19304 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		19578 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		19604 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		19701 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		19825 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		19875 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		19977 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		19980 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		20040 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		20157 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		20165 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		20217 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		20267 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		20283 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		20368 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		20419 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		20444 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		20520 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		20538 => STD_LOGIC_VECTOR(to_unsigned(182,8)),
		20542 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		20545 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		20738 => STD_LOGIC_VECTOR(to_unsigned(171,8)),
		20880 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		20918 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		20948 => STD_LOGIC_VECTOR(to_unsigned(77,8)),
		20981 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		21049 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		21052 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		21063 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		21111 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		21193 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		21301 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		21314 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		21325 => STD_LOGIC_VECTOR(to_unsigned(157,8)),
		21368 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		21388 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		21898 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		22054 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		22176 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		22245 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		22278 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		22286 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		22288 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		22311 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		22324 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		22490 => STD_LOGIC_VECTOR(to_unsigned(227,8)),
		22601 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		22657 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		22670 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		22688 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		22701 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		22904 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		22929 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		22965 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		23017 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		23086 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		23102 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		23186 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		23263 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		23281 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		23454 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		23567 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		23629 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		23647 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		23652 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		23692 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		23716 => STD_LOGIC_VECTOR(to_unsigned(134,8)),
		23832 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		24107 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		24138 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		24162 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		24233 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		24381 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		24429 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		24431 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		24451 => STD_LOGIC_VECTOR(to_unsigned(71,8)),
		24526 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		24609 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		24613 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		24617 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		24669 => STD_LOGIC_VECTOR(to_unsigned(94,8)),
		24733 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		24776 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		24898 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		25019 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		25064 => STD_LOGIC_VECTOR(to_unsigned(119,8)),
		25074 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		25108 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		25216 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		25268 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		25310 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		25449 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		25591 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		25600 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		25645 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		25673 => STD_LOGIC_VECTOR(to_unsigned(87,8)),
		25740 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		25791 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		25897 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		25908 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		25952 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		26051 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		26066 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		26161 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		26191 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		26244 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		26370 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		26435 => STD_LOGIC_VECTOR(to_unsigned(9,8)),
		26475 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		26724 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		26782 => STD_LOGIC_VECTOR(to_unsigned(140,8)),
		26838 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		26887 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		26902 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		26913 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		26915 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		26923 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		26929 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		26949 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		26985 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		27113 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		27161 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		27218 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		27276 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		27469 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		27523 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		27529 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		27548 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		27683 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		27792 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		27808 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		27919 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		28024 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		28062 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		28282 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		28437 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		28464 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		28562 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		28580 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		28634 => STD_LOGIC_VECTOR(to_unsigned(35,8)),
		28668 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		28755 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		28757 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		28765 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		28935 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		28944 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		29023 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		29051 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		29067 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		29101 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		29188 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		29240 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		29283 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		29292 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		29300 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		29315 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		29488 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		29493 => STD_LOGIC_VECTOR(to_unsigned(89,8)),
		29517 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		29535 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		29718 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		29750 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		29784 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		29893 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		29968 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		29974 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		29996 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		30130 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		30276 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		30371 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		30388 => STD_LOGIC_VECTOR(to_unsigned(5,8)),
		30407 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		30452 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		30556 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		30559 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		30561 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		30589 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		30753 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		30795 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		30805 => STD_LOGIC_VECTOR(to_unsigned(254,8)),
		30843 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		30952 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		30993 => STD_LOGIC_VECTOR(to_unsigned(42,8)),
		31033 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		31233 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		31240 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		31287 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		31298 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		31351 => STD_LOGIC_VECTOR(to_unsigned(176,8)),
		31479 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		31587 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		31619 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		31861 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		31881 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		31895 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		31916 => STD_LOGIC_VECTOR(to_unsigned(128,8)),
		31925 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		31938 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		32028 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		32066 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		32085 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		32187 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		32223 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		32305 => STD_LOGIC_VECTOR(to_unsigned(173,8)),
		32385 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		32412 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		32443 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		32457 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		32464 => STD_LOGIC_VECTOR(to_unsigned(124,8)),
		32620 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		32656 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		32686 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		32765 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		32915 => STD_LOGIC_VECTOR(to_unsigned(234,8)),
		32919 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		32999 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		33146 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		33476 => STD_LOGIC_VECTOR(to_unsigned(115,8)),
		33524 => STD_LOGIC_VECTOR(to_unsigned(195,8)),
		33570 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		33596 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		33618 => STD_LOGIC_VECTOR(to_unsigned(17,8)),
		33727 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		33759 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		33834 => STD_LOGIC_VECTOR(to_unsigned(211,8)),
		34022 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		34043 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		34072 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		34115 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		34206 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		34213 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		34317 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		34602 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		34659 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		34846 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		34859 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		34930 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		34983 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		35088 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		35124 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		35145 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		35325 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		35331 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		35381 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		35413 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		35431 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		35525 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		35627 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		35785 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		35862 => STD_LOGIC_VECTOR(to_unsigned(34,8)),
		36010 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		36016 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		36019 => STD_LOGIC_VECTOR(to_unsigned(144,8)),
		36063 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		36102 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		36159 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		36165 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		36219 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		36231 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		36316 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		36357 => STD_LOGIC_VECTOR(to_unsigned(230,8)),
		36397 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		36531 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		36604 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		36702 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		36705 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		36782 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		36844 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		36857 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		36947 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		37126 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		37132 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		37216 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		37386 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		37431 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		37476 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		37622 => STD_LOGIC_VECTOR(to_unsigned(50,8)),
		37664 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		37782 => STD_LOGIC_VECTOR(to_unsigned(160,8)),
		37819 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		37829 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		37830 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		37871 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		37882 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		37933 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		38062 => STD_LOGIC_VECTOR(to_unsigned(10,8)),
		38107 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		38141 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		38181 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		38195 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		38239 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		38441 => STD_LOGIC_VECTOR(to_unsigned(45,8)),
		38450 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		38575 => STD_LOGIC_VECTOR(to_unsigned(136,8)),
		38632 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		38715 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		38925 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		38929 => STD_LOGIC_VECTOR(to_unsigned(102,8)),
		38947 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		38968 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		39045 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		39167 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		39227 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		39284 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		39368 => STD_LOGIC_VECTOR(to_unsigned(247,8)),
		39426 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		39598 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		39638 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		39825 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		39989 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		40004 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		40016 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		40026 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		40109 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		40155 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		40283 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		40351 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		40470 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		40526 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		40677 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		40687 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		40713 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		41517 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		41546 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		41621 => STD_LOGIC_VECTOR(to_unsigned(67,8)),
		41889 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		41937 => STD_LOGIC_VECTOR(to_unsigned(59,8)),
		41938 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		41945 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		42035 => STD_LOGIC_VECTOR(to_unsigned(61,8)),
		42080 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		42104 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		42186 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		42195 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		42259 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		42404 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		42422 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		42423 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		42472 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		42600 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		42605 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		42951 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		43007 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		43040 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		43105 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		43169 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		43178 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		43250 => STD_LOGIC_VECTOR(to_unsigned(13,8)),
		43438 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		43604 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		43630 => STD_LOGIC_VECTOR(to_unsigned(250,8)),
		43705 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		43822 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		43839 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		43856 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		43937 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		43949 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		44065 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		44140 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		44196 => STD_LOGIC_VECTOR(to_unsigned(155,8)),
		44244 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		44306 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		44484 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		44574 => STD_LOGIC_VECTOR(to_unsigned(92,8)),
		44588 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		44702 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		44716 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		44723 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		44768 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		45087 => STD_LOGIC_VECTOR(to_unsigned(235,8)),
		45102 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		45111 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		45170 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		45237 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		45241 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		45258 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		45323 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		45404 => STD_LOGIC_VECTOR(to_unsigned(39,8)),
		45641 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		45660 => STD_LOGIC_VECTOR(to_unsigned(101,8)),
		45678 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		45705 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		45896 => STD_LOGIC_VECTOR(to_unsigned(20,8)),
		45909 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		46001 => STD_LOGIC_VECTOR(to_unsigned(204,8)),
		46083 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		46102 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		46196 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		46209 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		46245 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		46340 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		46382 => STD_LOGIC_VECTOR(to_unsigned(6,8)),
		46394 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		46458 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		46526 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		46589 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		46659 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		46719 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		46803 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		47026 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		47038 => STD_LOGIC_VECTOR(to_unsigned(133,8)),
		47101 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		47118 => STD_LOGIC_VECTOR(to_unsigned(201,8)),
		47143 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		47173 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		47225 => STD_LOGIC_VECTOR(to_unsigned(96,8)),
		47256 => STD_LOGIC_VECTOR(to_unsigned(229,8)),
		47421 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		47513 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		47523 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		47678 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		47830 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		47953 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		47987 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		48056 => STD_LOGIC_VECTOR(to_unsigned(158,8)),
		48225 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		48294 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		48336 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		48475 => STD_LOGIC_VECTOR(to_unsigned(82,8)),
		48534 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		48630 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		48631 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		48757 => STD_LOGIC_VECTOR(to_unsigned(154,8)),
		48814 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		48883 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		48891 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		48918 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		49082 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		49106 => STD_LOGIC_VECTOR(to_unsigned(28,8)),
		49132 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		49290 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		49536 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		49634 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		49670 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		49750 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		49785 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		49822 => STD_LOGIC_VECTOR(to_unsigned(207,8)),
		49935 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		49985 => STD_LOGIC_VECTOR(to_unsigned(72,8)),
		50173 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		50197 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		50254 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		50328 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		50373 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		50376 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		50410 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		50435 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		50438 => STD_LOGIC_VECTOR(to_unsigned(126,8)),
		50764 => STD_LOGIC_VECTOR(to_unsigned(83,8)),
		50824 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		50834 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		50903 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		50905 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		50910 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		50930 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		50953 => STD_LOGIC_VECTOR(to_unsigned(114,8)),
		51022 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		51040 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		51070 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		51078 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		51202 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		51266 => STD_LOGIC_VECTOR(to_unsigned(79,8)),
		51295 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		51314 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		51375 => STD_LOGIC_VECTOR(to_unsigned(248,8)),
		51444 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		51449 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		51485 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		51558 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		51579 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		51810 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		52012 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		52044 => STD_LOGIC_VECTOR(to_unsigned(107,8)),
		52078 => STD_LOGIC_VECTOR(to_unsigned(54,8)),
		52127 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		52319 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		52361 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		52362 => STD_LOGIC_VECTOR(to_unsigned(139,8)),
		52386 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		52419 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		52477 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		52557 => STD_LOGIC_VECTOR(to_unsigned(187,8)),
		52562 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		52578 => STD_LOGIC_VECTOR(to_unsigned(237,8)),
		52665 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		52745 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		52927 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		52945 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		52949 => STD_LOGIC_VECTOR(to_unsigned(209,8)),
		53016 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		53026 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		53066 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		53137 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		53208 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		53218 => STD_LOGIC_VECTOR(to_unsigned(131,8)),
		53236 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		53264 => STD_LOGIC_VECTOR(to_unsigned(110,8)),
		53307 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		53329 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		53391 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		53414 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		53578 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		53615 => STD_LOGIC_VECTOR(to_unsigned(129,8)),
		53687 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		53695 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		53704 => STD_LOGIC_VECTOR(to_unsigned(84,8)),
		53729 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		53785 => STD_LOGIC_VECTOR(to_unsigned(104,8)),
		53828 => STD_LOGIC_VECTOR(to_unsigned(146,8)),
		53845 => STD_LOGIC_VECTOR(to_unsigned(143,8)),
		53862 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		53881 => STD_LOGIC_VECTOR(to_unsigned(120,8)),
		53978 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		54116 => STD_LOGIC_VECTOR(to_unsigned(27,8)),
		54121 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		54133 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		54199 => STD_LOGIC_VECTOR(to_unsigned(196,8)),
		54241 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		54361 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		54364 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		54385 => STD_LOGIC_VECTOR(to_unsigned(52,8)),
		54398 => STD_LOGIC_VECTOR(to_unsigned(55,8)),
		54421 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		54526 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		54686 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		54703 => STD_LOGIC_VECTOR(to_unsigned(64,8)),
		54927 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		54982 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		55001 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		55034 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		55186 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		55226 => STD_LOGIC_VECTOR(to_unsigned(172,8)),
		55241 => STD_LOGIC_VECTOR(to_unsigned(69,8)),
		55282 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		55365 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		55543 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		55646 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		55834 => STD_LOGIC_VECTOR(to_unsigned(188,8)),
		55906 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		56006 => STD_LOGIC_VECTOR(to_unsigned(81,8)),
		56012 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		56046 => STD_LOGIC_VECTOR(to_unsigned(202,8)),
		56108 => STD_LOGIC_VECTOR(to_unsigned(58,8)),
		56134 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		56357 => STD_LOGIC_VECTOR(to_unsigned(98,8)),
		56441 => STD_LOGIC_VECTOR(to_unsigned(199,8)),
		56464 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		56507 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		56546 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		56551 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		56766 => STD_LOGIC_VECTOR(to_unsigned(49,8)),
		56820 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		56855 => STD_LOGIC_VECTOR(to_unsigned(132,8)),
		56866 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		56906 => STD_LOGIC_VECTOR(to_unsigned(112,8)),
		56925 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		57028 => STD_LOGIC_VECTOR(to_unsigned(36,8)),
		57106 => STD_LOGIC_VECTOR(to_unsigned(73,8)),
		57185 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		57280 => STD_LOGIC_VECTOR(to_unsigned(233,8)),
		57287 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		57419 => STD_LOGIC_VECTOR(to_unsigned(169,8)),
		57447 => STD_LOGIC_VECTOR(to_unsigned(25,8)),
		57515 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		57527 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		57544 => STD_LOGIC_VECTOR(to_unsigned(23,8)),
		57628 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		57781 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		57789 => STD_LOGIC_VECTOR(to_unsigned(70,8)),
		57806 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		57874 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		57883 => STD_LOGIC_VECTOR(to_unsigned(48,8)),
		57884 => STD_LOGIC_VECTOR(to_unsigned(76,8)),
		57899 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		57913 => STD_LOGIC_VECTOR(to_unsigned(29,8)),
		57946 => STD_LOGIC_VECTOR(to_unsigned(8,8)),
		58041 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		58078 => STD_LOGIC_VECTOR(to_unsigned(109,8)),
		58166 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		58197 => STD_LOGIC_VECTOR(to_unsigned(80,8)),
		58237 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		58242 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		58259 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		58268 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		58342 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		58364 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		58481 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		58485 => STD_LOGIC_VECTOR(to_unsigned(198,8)),
		58491 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		58535 => STD_LOGIC_VECTOR(to_unsigned(167,8)),
		58732 => STD_LOGIC_VECTOR(to_unsigned(63,8)),
		58969 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		59024 => STD_LOGIC_VECTOR(to_unsigned(252,8)),
		59037 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		59092 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		59189 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		59224 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		59332 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		59363 => STD_LOGIC_VECTOR(to_unsigned(74,8)),
		59461 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		59474 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		59482 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		59575 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		59656 => STD_LOGIC_VECTOR(to_unsigned(7,8)),
		59682 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		59775 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		59854 => STD_LOGIC_VECTOR(to_unsigned(66,8)),
		59856 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		59907 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		59917 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		59928 => STD_LOGIC_VECTOR(to_unsigned(103,8)),
		60095 => STD_LOGIC_VECTOR(to_unsigned(106,8)),
		60175 => STD_LOGIC_VECTOR(to_unsigned(161,8)),
		60184 => STD_LOGIC_VECTOR(to_unsigned(240,8)),
		60323 => STD_LOGIC_VECTOR(to_unsigned(153,8)),
		60340 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		60427 => STD_LOGIC_VECTOR(to_unsigned(193,8)),
		60525 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		60545 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		60642 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		60656 => STD_LOGIC_VECTOR(to_unsigned(88,8)),
		60674 => STD_LOGIC_VECTOR(to_unsigned(183,8)),
		60682 => STD_LOGIC_VECTOR(to_unsigned(2,8)),
		60701 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		60741 => STD_LOGIC_VECTOR(to_unsigned(135,8)),
		60749 => STD_LOGIC_VECTOR(to_unsigned(32,8)),
		60779 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		60937 => STD_LOGIC_VECTOR(to_unsigned(60,8)),
		60973 => STD_LOGIC_VECTOR(to_unsigned(41,8)),
		60983 => STD_LOGIC_VECTOR(to_unsigned(190,8)),
		61004 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		61042 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		61148 => STD_LOGIC_VECTOR(to_unsigned(170,8)),
		61172 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		61223 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		61346 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		61507 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		61658 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		61684 => STD_LOGIC_VECTOR(to_unsigned(178,8)),
		61752 => STD_LOGIC_VECTOR(to_unsigned(164,8)),
		61807 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		61826 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		61832 => STD_LOGIC_VECTOR(to_unsigned(255,8)),
		61854 => STD_LOGIC_VECTOR(to_unsigned(19,8)),
		61920 => STD_LOGIC_VECTOR(to_unsigned(150,8)),
		61925 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		61993 => STD_LOGIC_VECTOR(to_unsigned(226,8)),
		62079 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		62347 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		62399 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		62490 => STD_LOGIC_VECTOR(to_unsigned(116,8)),
		62495 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		62732 => STD_LOGIC_VECTOR(to_unsigned(85,8)),
		62794 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		62893 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		62910 => STD_LOGIC_VECTOR(to_unsigned(206,8)),
		62972 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		63043 => STD_LOGIC_VECTOR(to_unsigned(179,8)),
		63172 => STD_LOGIC_VECTOR(to_unsigned(177,8)),
		63183 => STD_LOGIC_VECTOR(to_unsigned(148,8)),
		63184 => STD_LOGIC_VECTOR(to_unsigned(21,8)),
		63230 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		63271 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		63301 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		63310 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		63363 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		63375 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		63386 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		63462 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		63532 => STD_LOGIC_VECTOR(to_unsigned(4,8)),
		63731 => STD_LOGIC_VECTOR(to_unsigned(225,8)),
		63769 => STD_LOGIC_VECTOR(to_unsigned(141,8)),
		63935 => STD_LOGIC_VECTOR(to_unsigned(203,8)),
		63967 => STD_LOGIC_VECTOR(to_unsigned(11,8)),
		64071 => STD_LOGIC_VECTOR(to_unsigned(44,8)),
		64183 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		64184 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		64217 => STD_LOGIC_VECTOR(to_unsigned(253,8)),
		64447 => STD_LOGIC_VECTOR(to_unsigned(117,8)),
		64465 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		64515 => STD_LOGIC_VECTOR(to_unsigned(118,8)),
		64560 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		64561 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		64578 => STD_LOGIC_VECTOR(to_unsigned(51,8)),
		64624 => STD_LOGIC_VECTOR(to_unsigned(33,8)),
		64658 => STD_LOGIC_VECTOR(to_unsigned(99,8)),
		64819 => STD_LOGIC_VECTOR(to_unsigned(212,8)),
		64903 => STD_LOGIC_VECTOR(to_unsigned(113,8)),
		65010 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		65054 => STD_LOGIC_VECTOR(to_unsigned(142,8)),
		65090 => STD_LOGIC_VECTOR(to_unsigned(127,8)),
		65140 => STD_LOGIC_VECTOR(to_unsigned(214,8)),
		65149 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		65530 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		65535 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		others => (others => '0')
	);

	COMPONENT project_reti_logiche IS
		PORT (
			i_clk : IN STD_LOGIC;
			i_rst : IN STD_LOGIC;
			i_start : IN STD_LOGIC;
			i_w : IN STD_LOGIC;

			o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_done : OUT STD_LOGIC;

			o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_mem_we : OUT STD_LOGIC;
			o_mem_en : OUT STD_LOGIC
		);
	END COMPONENT project_reti_logiche;

BEGIN
	UUT : project_reti_logiche
	PORT MAP(
		i_clk => tb_clk,
		i_start => tb_start,
		i_rst => tb_rst,
		i_w => tb_w,

		o_z0 => tb_z0,
		o_z1 => tb_z1,
		o_z2 => tb_z2,
		o_z3 => tb_z3,
		o_done => tb_done,

		o_mem_addr => mem_address,
		o_mem_en => enable_wire,
		o_mem_we => mem_we,
		i_mem_data => mem_o_data
	);


	-- Process for the clock generation
	CLK_GEN : PROCESS IS
	BEGIN
		WAIT FOR CLOCK_PERIOD/2;
		tb_clk <= NOT tb_clk;
	END PROCESS CLK_GEN;


	-- Process related to the memory
	MEM : PROCESS (tb_clk)
	BEGIN
		IF tb_clk'event AND tb_clk = '1' THEN
			IF enable_wire = '1' THEN
				IF mem_we = '1' THEN
					RAM(conv_integer(mem_address)) <= mem_i_data;
					mem_o_data <= mem_i_data AFTER 1 ns;
				ELSE
					mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns;
				END IF;
			END IF;
		END IF;
	END PROCESS;

	-- This process provides the correct scenario on the signal controlled by the TB
	createScenario : PROCESS (tb_clk)
	BEGIN
		IF tb_clk'event AND tb_clk = '0' THEN
			tb_rst <= scenario_rst(0);
			tb_w <= scenario_w(0);
			tb_start <= scenario_start(0);
			scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
			scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
			scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
		END IF;
	END PROCESS;

	-- Process without sensitivity list designed to test the actual component.
	testRoutine : PROCESS IS
	BEGIN
		FOR i IN 0 TO N_EVENTS - 1 LOOP
			mem_i_data <= "00000000";
			IF do_reset(i) = '1' THEN
				WAIT UNTIL tb_rst = '1';
				WAIT UNTIL tb_rst = '0';
				ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure;
				ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure;
				ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
				ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
				ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset done != 0 )" severity failure;
				ASSERT enable_wire = '0' REPORT "TEST FALLITO (postreset enable_wire != 0 )" severity warning;
				ASSERT mem_we = '0' REPORT "(mem_we != 0 )" severity failure;
			END IF;

			WAIT UNTIL tb_start = '1';
			ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure;
			ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure;
			ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
			ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure;
			ASSERT tb_done = '0' REPORT "TEST FALLITO (poststart done != 0 )" severity failure;
			ASSERT enable_wire = '0' REPORT "TEST FALLITO (poststart enable_wire != 0 )" severity warning;
			ASSERT mem_we = '0' REPORT "(mem_we != 0 )" severity failure;
			WAIT UNTIL tb_done = '1';
			--WAIT UNTIL rising_edge(tb_clk);
			WAIT FOR CLOCK_PERIOD/2;
			ASSERT tb_z0 = std_logic_vector(to_unsigned(registers_check(i, 0), 8))	REPORT "TEST FALLITO (Z0 ---) found " & integer'image(to_integer(unsigned(tb_z0))) & " Expected " & integer'image(registers_check(i, 0)) severity failure;
			ASSERT tb_z1 = std_logic_vector(to_unsigned(registers_check(i, 1), 8))	REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z1))) & " Expected " & integer'image(registers_check(i, 1)) severity failure;
			ASSERT tb_z2 = std_logic_vector(to_unsigned(registers_check(i, 2), 8))	REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z2))) & " Expected " & integer'image(registers_check(i, 2)) severity failure;
			ASSERT tb_z3 = std_logic_vector(to_unsigned(registers_check(i, 3), 8))	REPORT "TEST FALLITO (Z3 ---) found " & integer'image(to_integer(unsigned(tb_z3))) & " Expected " & integer'image(registers_check(i, 3)) severity failure;
			ASSERT tb_done = '1' REPORT "TEST FALLITO (done = 0 )" severity failure;
			WAIT FOR CLOCK_PERIOD/2 + 10 ns;
			ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure;
			ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure;
			ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
			ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure;
			ASSERT tb_done = '0' REPORT "TEST FALLITO (postdone done != 0 )" severity failure;
			ASSERT enable_wire = '0' REPORT "(postdone enable_wire != 0 )" severity warning;
			ASSERT mem_we = '0' REPORT "TEST FALLITO (mem_we != 0 )" severity failure;
		END LOOP;
		wait FOR CLOCK_PERIOD * 2;
		REPORT "SUCCESS";
		finish;
	END PROCESS testRoutine;

END randomtb;

