
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;
USE std.env.finish;

ENTITY random_tb IS
END random_tb;

ARCHITECTURE randomtb OF random_tb IS
	CONSTANT CLOCK_PERIOD : TIME := 100 ns;
	SIGNAL tb_done : STD_LOGIC;
	SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
	SIGNAL tb_rst : STD_LOGIC := '0';
	SIGNAL tb_start : STD_LOGIC := '0';
	SIGNAL tb_clk : STD_LOGIC := '0';
	SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL enable_wire : STD_LOGIC;
	SIGNAL mem_we : STD_LOGIC;
	SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL tb_w : STD_LOGIC;

	CONSTANT SCENARIOLENGTH : INTEGER := 4071;
	CONSTANT N_EVENTS : INTEGER := 100;
	SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)		:= "010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000010000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
	SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)	:= "000011111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111000000000000000000000111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111100000000000000000000000111111111111111000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000111111111111111100000000000000000000000111111111111111111000000000000000000001000001111111111111111110000000000000000000000000011111111111111111000000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111110000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111110000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000001111111111111111000000000000000000000000111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000001111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000000001111111111111111110000000000000000000001111111111111111110000000000000000000000111111111111111111000000000000000000000011111111111111100000000000000000000000001111111111111111000000000000000000000011111111111111111000000000000000000000000011111111111111111000000000000000000000001111111111111111110000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000001111111111111111110000000000000000000000000111111111111111110000000000000000000000000111111111111111000000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000111111111111111100000000000000000000100111111111111111111000000000000000000000111111111111111111000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000011111111111111111000000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000100011111111111111111000000000000000000000000011111111111111111100000000000000000000000001111111111111111110000000000000000000000000111111111111111111000000000000000000000011111111111111111000000000000000000000111111111111111111000000000000000000000000011111111111111111100000000000000000000000011111111111111111100000000000000000000000111111111111111110000000000000000000000000111111111111111111000000000000000000000111111111111111111000000000000000000000011111111111111111100000000000000000000000111111111111111100000000000000000000011111111111111111100000000000000000000";
	SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)		:= "011101110100011011001110010010110001110101001111011011110101110111100001101011110110011011111001110111010001001100001011101110000111111110010101101110010010111110000100111100010011100001110111101100000110110011010011110100100011010000111101011000100010100000100001101100000111100111011101110011011101111001101101001000101110110101111010101011101000001100000001011111010111111011011001110100000001101101000010000011001001110011111001001010100100111010000011111111101100011101100010000100100010111100111111110111010011100100001010010110110001100001111010000000000011001100110010110100110110110000111010011001100110011001111001101101010101101000011110110101000010101011011001110110100011111111100100100100001010001001011000011000100110101110111111000100111010111110100110100100010010110111100010010100011111110010010100011000010011001101000010011100101111010101110111001010000100011010100001010010001111111011110110000110101110110011001111001100011111000011001101011101100010011110100100100000110100101101110011001011100110110000111111001001111100001011000001111000101000100111010011000111110111101101100100101111001000011110100001000001001000010001010110011100111111001101111010111001011011000100011010110001001010101100000100001011001010001001101000000011101100100110001010111111000111001001101000111101100011001000001010001111011001001101101010111110010011001101101011001100100100100110101001010010010100001111111001110011001101001100110000101001001110101101001010011010111011000010011001100100101011010110000010111101110000000011011111001001111001001000110011010001000011111011001010010100110110010010110000101110010011001000110000001001001000001011110111000110001101110001110101111011111010110100011111111101110100111011001100011111110000000011011100101001000000010100001100110100001001110111101001110110001100011001010111010010111101111011101111011011101111111100010000110100001111100101111000011100101100010100001101000010001000110000000011100100111110101100111110101100100010110111001001010010000110101110111010010101011001000101001000011101010110010110111100001110001011110100101001010101000011001100000111111011011000011100001100010100111011100110100010010110011111011000011101100011110111001011011100010001111110100100111110011101010110111100111101010101010011011100010111100111000101010011010111000001100111001110100100010111010101011111101000000100010011110110111011110100001000001001111111110101010010010111101011110111111100010100001111010001000111000011000010000010010010110001100111001111110010110010101101000010001011100100111011001010011011101010100101111100011001100110010101110100110011001001011000010110111110100000001001000001010000001010100101000101101101111110101001001111000000000010100011111011100011110010100000000100010011010111011101111110111001011001101101111101000010100110111101111010001100100100100001100000011101010100111100100010110010011101110110101001100011001000011010110100100001111111100111101011001101101111000010100100100001000101111000111011000000000010100110000001011101000111100010100001010110111110101011000011100101001101010010110010000010010100100100011110011000010001110111010010111011101101101001011001110001100011110111000010011001011011000101010010110010111011100010000011111010000011011001001001011000111000000100001001001111001100010110110011010010101110111000111100000000110001000010100000111011000101000110010110000110011110000111100111110000011001111101101001100011111011010010111011010111100101011010101010101010001011001101011101101001001011110011010000110111001001001010110101110101110110101010101101110010000011010000000010101001010100010111001101111110000010100011001100101101001010110101011011101011101000011110100101001101101010011101011001001100110110111010001110111000111111111100001010101101111001000011001111011100011001110010111111101101111110001011100111011110011000011000110110101100111001101001001010011001111000000010110000011100100101010011000101111110000110101100000100010001111000100010101010100010000101101111011010010000100110100100011001011101111001101100110001011111001101001110001001101101101";

	TYPE registers IS ARRAY (0 TO N_EVENTS - 1, 0 TO 3) OF INTEGER;
	SIGNAL registers_check : registers := (
		(0,105,0,0),(0,166,0,0),(0,166,0,217),(123,166,0,217),(123,166,130,217),(123,56,130,217),(0,0,0,100),(0,151,0,100),(0,93,0,100),(0,93,0,221),(0,222,0,221),(0,222,0,200),(0,191,0,200),(238,0,0,0),(238,0,12,0),(238,0,159,0),(238,0,159,231),(238,0,159,224),(220,0,159,224),(220,0,189,224),(220,0,189,152),(0,245,0,0),(0,0,86,0),(0,121,86,0),(0,223,0,0),(47,223,0,0),(47,223,0,122),(215,223,0,122),(26,223,0,122),(228,223,0,122),(218,223,0,122),(218,239,0,122),(97,239,0,122),(97,239,90,122),(97,46,90,122),(97,46,216,122),(97,46,244,122),(97,46,184,122),(97,46,147,122),(97,220,147,122),(186,220,147,122),(186,197,147,122),(186,197,147,165),(186,197,189,165),(0,0,0,14),(0,0,0,152),(236,0,0,152),(236,38,0,152),(0,0,0,210),(0,0,241,210),(0,0,1,210),(0,57,1,210),(0,57,1,53),(192,57,1,53),(192,57,185,53),(156,57,185,53),(162,57,185,53),(0,0,0,0),(138,0,0,0),(138,0,0,123),(138,243,0,123),(138,111,0,123),(138,111,47,123),(138,111,75,123),(138,111,175,123),(251,111,175,123),(0,0,168,0),(0,232,168,0),(0,232,168,181),(0,232,24,181),(0,239,24,181),(0,174,24,181),(0,0,0,208),(0,0,30,208),(0,0,219,208),(53,0,219,208),(194,0,219,208),(194,242,219,208),(91,242,219,208),(145,242,219,208),(65,242,219,208),(65,242,163,208),(65,242,78,208),(65,242,180,208),(65,249,180,208),(65,249,205,208),(0,0,0,40),(0,0,125,40),(0,0,210,40),(0,0,37,40),(0,0,130,40),(0,0,130,122),(0,213,130,122),(0,213,130,15),(0,68,130,15),(0,68,130,205),(0,68,220,205),(246,68,220,205),(246,68,22,205),(246,68,192,205)
	);

	SIGNAL do_reset : std_logic_vector(0 TO N_EVENTS - 1) := "1000001000000100000001101000000000000000000010001000000001000000001000001000000000000010000000000000";

	TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL RAM : ram_type := (
		241 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		310 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		1420 => STD_LOGIC_VECTOR(to_unsigned(111,8)),
		1614 => STD_LOGIC_VECTOR(to_unsigned(222,8)),
		3036 => STD_LOGIC_VECTOR(to_unsigned(184,8)),
		3252 => STD_LOGIC_VECTOR(to_unsigned(12,8)),
		3914 => STD_LOGIC_VECTOR(to_unsigned(57,8)),
		4417 => STD_LOGIC_VECTOR(to_unsigned(100,8)),
		4659 => STD_LOGIC_VECTOR(to_unsigned(147,8)),
		6047 => STD_LOGIC_VECTOR(to_unsigned(191,8)),
		6125 => STD_LOGIC_VECTOR(to_unsigned(221,8)),
		6405 => STD_LOGIC_VECTOR(to_unsigned(97,8)),
		6558 => STD_LOGIC_VECTOR(to_unsigned(159,8)),
		6724 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		6726 => STD_LOGIC_VECTOR(to_unsigned(22,8)),
		7804 => STD_LOGIC_VECTOR(to_unsigned(180,8)),
		8633 => STD_LOGIC_VECTOR(to_unsigned(40,8)),
		8680 => STD_LOGIC_VECTOR(to_unsigned(243,8)),
		9211 => STD_LOGIC_VECTOR(to_unsigned(86,8)),
		9825 => STD_LOGIC_VECTOR(to_unsigned(216,8)),
		10261 => STD_LOGIC_VECTOR(to_unsigned(251,8)),
		12186 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		13855 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		14019 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		14917 => STD_LOGIC_VECTOR(to_unsigned(0,8)),
		15675 => STD_LOGIC_VECTOR(to_unsigned(14,8)),
		16884 => STD_LOGIC_VECTOR(to_unsigned(145,8)),
		17218 => STD_LOGIC_VECTOR(to_unsigned(38,8)),
		17767 => STD_LOGIC_VECTOR(to_unsigned(26,8)),
		18134 => STD_LOGIC_VECTOR(to_unsigned(68,8)),
		18675 => STD_LOGIC_VECTOR(to_unsigned(194,8)),
		19053 => STD_LOGIC_VECTOR(to_unsigned(130,8)),
		19211 => STD_LOGIC_VECTOR(to_unsigned(175,8)),
		19638 => STD_LOGIC_VECTOR(to_unsigned(91,8)),
		19831 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		20258 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		21828 => STD_LOGIC_VECTOR(to_unsigned(246,8)),
		23320 => STD_LOGIC_VECTOR(to_unsigned(238,8)),
		26748 => STD_LOGIC_VECTOR(to_unsigned(236,8)),
		26774 => STD_LOGIC_VECTOR(to_unsigned(192,8)),
		26841 => STD_LOGIC_VECTOR(to_unsigned(105,8)),
		27568 => STD_LOGIC_VECTOR(to_unsigned(244,8)),
		28302 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		29338 => STD_LOGIC_VECTOR(to_unsigned(53,8)),
		29404 => STD_LOGIC_VECTOR(to_unsigned(185,8)),
		30453 => STD_LOGIC_VECTOR(to_unsigned(166,8)),
		30542 => STD_LOGIC_VECTOR(to_unsigned(165,8)),
		31419 => STD_LOGIC_VECTOR(to_unsigned(245,8)),
		31982 => STD_LOGIC_VECTOR(to_unsigned(217,8)),
		32661 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		32944 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		33713 => STD_LOGIC_VECTOR(to_unsigned(78,8)),
		33884 => STD_LOGIC_VECTOR(to_unsigned(47,8)),
		34196 => STD_LOGIC_VECTOR(to_unsigned(218,8)),
		35309 => STD_LOGIC_VECTOR(to_unsigned(138,8)),
		35367 => STD_LOGIC_VECTOR(to_unsigned(122,8)),
		35580 => STD_LOGIC_VECTOR(to_unsigned(239,8)),
		35849 => STD_LOGIC_VECTOR(to_unsigned(186,8)),
		35974 => STD_LOGIC_VECTOR(to_unsigned(174,8)),
		36628 => STD_LOGIC_VECTOR(to_unsigned(219,8)),
		37079 => STD_LOGIC_VECTOR(to_unsigned(241,8)),
		37098 => STD_LOGIC_VECTOR(to_unsigned(1,8)),
		37824 => STD_LOGIC_VECTOR(to_unsigned(168,8)),
		38364 => STD_LOGIC_VECTOR(to_unsigned(163,8)),
		38800 => STD_LOGIC_VECTOR(to_unsigned(215,8)),
		38854 => STD_LOGIC_VECTOR(to_unsigned(75,8)),
		41215 => STD_LOGIC_VECTOR(to_unsigned(200,8)),
		41702 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		43187 => STD_LOGIC_VECTOR(to_unsigned(205,8)),
		43337 => STD_LOGIC_VECTOR(to_unsigned(46,8)),
		43740 => STD_LOGIC_VECTOR(to_unsigned(125,8)),
		44251 => STD_LOGIC_VECTOR(to_unsigned(208,8)),
		44282 => STD_LOGIC_VECTOR(to_unsigned(210,8)),
		44885 => STD_LOGIC_VECTOR(to_unsigned(93,8)),
		45903 => STD_LOGIC_VECTOR(to_unsigned(56,8)),
		46627 => STD_LOGIC_VECTOR(to_unsigned(228,8)),
		47339 => STD_LOGIC_VECTOR(to_unsigned(197,8)),
		47462 => STD_LOGIC_VECTOR(to_unsigned(181,8)),
		48262 => STD_LOGIC_VECTOR(to_unsigned(213,8)),
		48354 => STD_LOGIC_VECTOR(to_unsigned(162,8)),
		48716 => STD_LOGIC_VECTOR(to_unsigned(90,8)),
		53941 => STD_LOGIC_VECTOR(to_unsigned(37,8)),
		55941 => STD_LOGIC_VECTOR(to_unsigned(231,8)),
		56139 => STD_LOGIC_VECTOR(to_unsigned(242,8)),
		56541 => STD_LOGIC_VECTOR(to_unsigned(151,8)),
		57071 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		57410 => STD_LOGIC_VECTOR(to_unsigned(65,8)),
		58531 => STD_LOGIC_VECTOR(to_unsigned(152,8)),
		58624 => STD_LOGIC_VECTOR(to_unsigned(232,8)),
		58656 => STD_LOGIC_VECTOR(to_unsigned(189,8)),
		58942 => STD_LOGIC_VECTOR(to_unsigned(121,8)),
		59680 => STD_LOGIC_VECTOR(to_unsigned(223,8)),
		60126 => STD_LOGIC_VECTOR(to_unsigned(156,8)),
		61912 => STD_LOGIC_VECTOR(to_unsigned(30,8)),
		62564 => STD_LOGIC_VECTOR(to_unsigned(24,8)),
		63127 => STD_LOGIC_VECTOR(to_unsigned(249,8)),
		63228 => STD_LOGIC_VECTOR(to_unsigned(15,8)),
		64565 => STD_LOGIC_VECTOR(to_unsigned(220,8)),
		65097 => STD_LOGIC_VECTOR(to_unsigned(224,8)),
		65193 => STD_LOGIC_VECTOR(to_unsigned(123,8)),
		others => (others => '0')
	);

	COMPONENT project_reti_logiche IS
		PORT (
			i_clk : IN STD_LOGIC;
			i_rst : IN STD_LOGIC;
			i_start : IN STD_LOGIC;
			i_w : IN STD_LOGIC;

			o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_done : OUT STD_LOGIC;

			o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
			i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			o_mem_we : OUT STD_LOGIC;
			o_mem_en : OUT STD_LOGIC
		);
	END COMPONENT project_reti_logiche;

BEGIN
	UUT : project_reti_logiche
	PORT MAP(
		i_clk => tb_clk,
		i_start => tb_start,
		i_rst => tb_rst,
		i_w => tb_w,

		o_z0 => tb_z0,
		o_z1 => tb_z1,
		o_z2 => tb_z2,
		o_z3 => tb_z3,
		o_done => tb_done,

		o_mem_addr => mem_address,
		o_mem_en => enable_wire,
		o_mem_we => mem_we,
		i_mem_data => mem_o_data
	);


	-- Process for the clock generation
	CLK_GEN : PROCESS IS
	BEGIN
		WAIT FOR CLOCK_PERIOD/2;
		tb_clk <= NOT tb_clk;
	END PROCESS CLK_GEN;


	-- Process related to the memory
	MEM : PROCESS (tb_clk)
	BEGIN
		IF tb_clk'event AND tb_clk = '1' THEN
			IF enable_wire = '1' THEN
				IF mem_we = '1' THEN
					RAM(conv_integer(mem_address)) <= mem_i_data;
					mem_o_data <= mem_i_data AFTER 1 ns;
				ELSE
					mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns;
				END IF;
			END IF;
		END IF;
	END PROCESS;

	-- This process provides the correct scenario on the signal controlled by the TB
	createScenario : PROCESS (tb_clk)
	BEGIN
		IF tb_clk'event AND tb_clk = '0' THEN
			tb_rst <= scenario_rst(0);
			tb_w <= scenario_w(0);
			tb_start <= scenario_start(0);
			scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
			scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
			scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
		END IF;
	END PROCESS;

	-- Process without sensitivity list designed to test the actual component.
	testRoutine : PROCESS IS
	BEGIN
		FOR i IN 0 TO N_EVENTS - 1 LOOP
			mem_i_data <= "00000000";
			IF do_reset(i) = '1' THEN
				WAIT UNTIL tb_rst = '1';
				WAIT UNTIL tb_rst = '0';
				ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure;
				ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure;
				ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
				ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postreset Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
				ASSERT tb_done = '0' REPORT "TEST FALLITO (postreset done != 0 )" severity failure;
				ASSERT enable_wire = '0' REPORT "TEST FALLITO (postreset enable_wire != 0 )" severity warning;
				ASSERT mem_we = '0' REPORT "(mem_we != 0 )" severity failure;
			END IF;

			WAIT UNTIL tb_start = '1';
			ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure;
			ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure;
			ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
			ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (poststart Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure;
			ASSERT tb_done = '0' REPORT "TEST FALLITO (poststart done != 0 )" severity failure;
			ASSERT enable_wire = '0' REPORT "TEST FALLITO (poststart enable_wire != 0 )" severity warning;
			ASSERT mem_we = '0' REPORT "(mem_we != 0 )" severity failure;
			WAIT UNTIL tb_done = '1';
			--WAIT UNTIL rising_edge(tb_clk);
			WAIT FOR CLOCK_PERIOD/2;
			ASSERT tb_z0 = std_logic_vector(to_unsigned(registers_check(i, 0), 8))	REPORT "TEST FALLITO (Z0 ---) found " & integer'image(to_integer(unsigned(tb_z0))) & " Expected " & integer'image(registers_check(i, 0)) severity failure;
			ASSERT tb_z1 = std_logic_vector(to_unsigned(registers_check(i, 1), 8))	REPORT "TEST FALLITO (Z1 ---) found " & integer'image(to_integer(unsigned(tb_z1))) & " Expected " & integer'image(registers_check(i, 1)) severity failure;
			ASSERT tb_z2 = std_logic_vector(to_unsigned(registers_check(i, 2), 8))	REPORT "TEST FALLITO (Z2 ---) found " & integer'image(to_integer(unsigned(tb_z2))) & " Expected " & integer'image(registers_check(i, 2)) severity failure;
			ASSERT tb_z3 = std_logic_vector(to_unsigned(registers_check(i, 3), 8))	REPORT "TEST FALLITO (Z3 ---) found " & integer'image(to_integer(unsigned(tb_z3))) & " Expected " & integer'image(registers_check(i, 3)) severity failure;
			ASSERT tb_done = '1' REPORT "TEST FALLITO (done = 0 )" severity failure;
			WAIT FOR CLOCK_PERIOD/2 + 10 ns;
			ASSERT tb_z0 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z0))) severity failure;
			ASSERT tb_z1 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z1))) severity failure;
			ASSERT tb_z2 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z2))) severity failure;
			ASSERT tb_z3 = "00000000" REPORT "TEST FALLITO (postdone Z0--Z3 != 0 ) found " & integer'image(to_integer(unsigned(tb_z3))) severity failure;
			ASSERT tb_done = '0' REPORT "TEST FALLITO (postdone done != 0 )" severity failure;
			ASSERT enable_wire = '0' REPORT "(postdone enable_wire != 0 )" severity warning;
			ASSERT mem_we = '0' REPORT "TEST FALLITO (mem_we != 0 )" severity failure;
		END LOOP;
		wait FOR CLOCK_PERIOD * 2;
		REPORT "SUCCESS";
		finish;
	END PROCESS testRoutine;

END randomtb;

