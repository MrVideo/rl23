-- Custom test bench 1
-- Tests for:
-- * 0 bit address
-- * Reset between runs

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.std_logic_unsigned.ALL;
USE std.textio.ALL;
USE std.env.finish;

ENTITY project_tb IS
END project_tb;

ARCHITECTURE projecttb OF project_tb IS
    CONSTANT CLOCK_PERIOD : TIME := 100 ns;
    SIGNAL tb_done : STD_LOGIC;
    SIGNAL mem_address : STD_LOGIC_VECTOR (15 DOWNTO 0) := (OTHERS => '0');
    SIGNAL tb_rst : STD_LOGIC := '0';
    SIGNAL tb_start : STD_LOGIC := '0';
    SIGNAL tb_clk : STD_LOGIC := '0';
    SIGNAL mem_o_data, mem_i_data : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL enable_wire : STD_LOGIC;
    SIGNAL mem_we : STD_LOGIC;
    SIGNAL tb_z0, tb_z1, tb_z2, tb_z3 : STD_LOGIC_VECTOR (7 DOWNTO 0);
    SIGNAL tb_w : STD_LOGIC;

    CONSTANT SCENARIOLENGTH : INTEGER := 428;
    SIGNAL scenario_rst : unsigned(0 TO SCENARIOLENGTH - 1)     := "00111111110000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000111111110000000000000000000000000000000000000000000000000001111111111111111000000000000000000000000111100000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001111111100000000000000000000000000000000001111111111000000000000000111111111111111111111111110000";
    SIGNAL scenario_start : unsigned(0 TO SCENARIOLENGTH - 1)   := "00000000000000000000000011000000000000000000000000000000000000000000000000000001100000000000000000000000000000000000000000011111111111111111100000000000000011111111000000000000001100000000000000000000000000110000000000000000111111111111111111000000000000000011111111000000000000000011111111110000000000000000111111111111111111000000000000000000000000000111111111111111111000000000000000111111110000000000000000000000000000000000";
    SIGNAL scenario_w : unsigned(0 TO SCENARIOLENGTH - 1)       := "00000000000000000000000010000000000000000000000000000000000000000000000000000000100000000000000000000000000000000000000000010111111111111111100000000000000000111110000011111111000100000000000000000000000000000000000000000000011111111111111111000000000000000010111111000000000000000011001100110000000000000000001111111111111111000000000000000000000000000101111111111111111000000000000000001111100000000000000000000000000000000000";
    -- Channel 2 -> MEM[1] -> 162
    -- Channel 1 -> MEM[2] -> 75

    TYPE ram_type IS ARRAY (65535 DOWNTO 0) OF STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL RAM : ram_type := (  0 => STD_LOGIC_VECTOR(to_unsigned(20, 8)), 
				1 => STD_LOGIC_VECTOR(to_unsigned(162, 8)), 
				2 => STD_LOGIC_VECTOR(to_unsigned(75, 8)), 
				3 => STD_LOGIC_VECTOR(to_unsigned(175, 8)), 
				6 => STD_LOGIC_VECTOR(to_unsigned(88, 8)), 
                51 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
				57 => STD_LOGIC_VECTOR(to_unsigned(18, 8)),
                62 => STD_LOGIC_VECTOR(to_unsigned(26, 8)),
                63 => STD_LOGIC_VECTOR(to_unsigned(9, 8)),  
				985 => STD_LOGIC_VECTOR(to_unsigned(456, 8)), 
				721 => STD_LOGIC_VECTOR(to_unsigned(98, 8)), 
				420 => STD_LOGIC_VECTOR(to_unsigned(420, 8)), 
				65535 => STD_LOGIC_VECTOR(to_unsigned(400, 8)), 
				1821 => STD_LOGIC_VECTOR(to_unsigned(697, 8)), 
				1312 => STD_LOGIC_VECTOR(to_unsigned(985, 8)), 
				7765 => STD_LOGIC_VECTOR(to_unsigned(894, 8)), 
				214 => STD_LOGIC_VECTOR(to_unsigned(59, 8)), 
				9 => STD_LOGIC_VECTOR(to_unsigned(654, 8)), 
				3059 => STD_LOGIC_VECTOR(to_unsigned(6, 8)), 
				69 => STD_LOGIC_VECTOR(to_unsigned(69, 8)), 
				 OTHERS => "00000000"-- (OTHERS => '0')
                            );

    COMPONENT project_reti_logiche IS
        PORT (
            i_clk : IN STD_LOGIC;
            i_rst : IN STD_LOGIC;
            i_start : IN STD_LOGIC;
            i_w : IN STD_LOGIC;

            o_z0 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z1 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z2 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_z3 : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_done : OUT STD_LOGIC;

            o_mem_addr : OUT STD_LOGIC_VECTOR(15 DOWNTO 0);
            i_mem_data : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
            o_mem_we : OUT STD_LOGIC;
            o_mem_en : OUT STD_LOGIC
        );
    END COMPONENT project_reti_logiche;

BEGIN
    UUT : project_reti_logiche
    PORT MAP(
        i_clk => tb_clk,
        i_start => tb_start,
        i_rst => tb_rst,
        i_w => tb_w,

        o_z0 => tb_z0,
        o_z1 => tb_z1,
        o_z2 => tb_z2,
        o_z3 => tb_z3,
        o_done => tb_done,

        o_mem_addr => mem_address,
        o_mem_en => enable_wire,
        o_mem_we => mem_we,
        i_mem_data => mem_o_data
    );


    -- Process for the clock generation
    CLK_GEN : PROCESS IS
    BEGIN
        WAIT FOR CLOCK_PERIOD/2;
        tb_clk <= NOT tb_clk;
    END PROCESS CLK_GEN;


    -- Process related to the memory
    MEM : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '1' THEN
            IF enable_wire = '1' THEN
                IF mem_we = '1' THEN
                    RAM(conv_integer(mem_address)) <= mem_i_data;
                    mem_o_data <= mem_i_data AFTER 1 ns;
                ELSE
                    mem_o_data <= RAM(conv_integer(mem_address)) AFTER 1 ns; 
                END IF;
            END IF;
        END IF;
    END PROCESS;

    -- This process provides the correct scenario on the signal controlled by the TB
    createScenario : PROCESS (tb_clk)
    BEGIN
        IF tb_clk'event AND tb_clk = '0' THEN
            tb_rst <= scenario_rst(0);
            tb_w <= scenario_w(0);
            tb_start <= scenario_start(0);
            scenario_rst <= scenario_rst(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_w <= scenario_w(1 TO SCENARIOLENGTH - 1) & '0';
            scenario_start <= scenario_start(1 TO SCENARIOLENGTH - 1) & '0';
        END IF;
    END PROCESS;

    -- Process without sensitivity list designed to test the actual component.
    testRoutine : PROCESS IS
    BEGIN
        mem_i_data <= "00000000";

        -- FIRST TEST
        
        -- First reset
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z3))) severity failure;
        
        -- First run
        WAIT UNTIL tb_start = '1';
        ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        
        WAIT UNTIL tb_done = '1';
        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
        ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
        ASSERT tb_z2 = std_logic_vector(to_unsigned(20, 8)) REPORT "Failed: Z0 was not 0x14" severity failure;
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
        WAIT UNTIL tb_done = '0';   
        
        -- Second reset
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z3))) severity failure;
        
        -- Second run
        WAIT UNTIL tb_start = '1';
        ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        
        WAIT UNTIL tb_done = '1';
        ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
        ASSERT tb_z1 = std_logic_vector(to_unsigned(20, 8)) REPORT "Failed: Z0 was not 0x14" severity failure;
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
        WAIT UNTIL tb_done = '0';   

        -- SECOND TEST

         -- First reset
         WAIT UNTIL tb_rst = '1';
         WAIT UNTIL tb_rst = '0';
         ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
         ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
         ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
         ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z3))) severity failure;
         
         -- First run
         WAIT UNTIL tb_start = '1';
         ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
         ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
         ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
         ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
         
         WAIT UNTIL tb_done = '1';
         ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
         ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
         ASSERT tb_z2 = std_logic_vector(to_unsigned(400, 8)) REPORT "Failed: Z0 was not 0x190" severity failure;
         ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
         WAIT UNTIL tb_done = '0';   
         
         -- Second run
         WAIT UNTIL tb_start = '1';
         ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
         ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
         ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
         ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure;
         
         -- Interruption by reset signal
         WAIT UNTIL tb_rst = '1';
         WAIT UNTIL tb_rst = '0';
         ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
         ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
         ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
         ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z3))) severity failure;
         
         -- Thrid run run
         WAIT UNTIL tb_start = '1';
         ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
         ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
         ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
         ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
         
         WAIT UNTIL tb_done = '1';
         ASSERT tb_z0 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
         ASSERT tb_z1 = std_logic_vector(to_unsigned(20, 8)) REPORT "Failed: Z0 was not 0x14" severity failure;
         ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
         ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z0 was not 0"  severity failure;
         WAIT UNTIL tb_done = '0';   
        
        -- THIRD TEST

        -- Reset
        WAIT UNTIL tb_rst = '1';
        WAIT UNTIL tb_rst = '0';
        ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z3))) severity failure;
        
        -- First run
        WAIT UNTIL tb_start = '1';
        ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        
        WAIT UNTIL tb_done = '1';
        ASSERT tb_z0 = std_logic_vector(to_unsigned(20, 8)) REPORT "Failed: Z0 was not 0x14" severity failure;
        ASSERT tb_z1 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z1 was not 0"    severity failure;
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z2 was not 0"    severity failure;
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))  REPORT "Failed: Z3 was not 0"    severity failure;
        WAIT UNTIL tb_done = '0';
        WAIT FOR CLOCK_PERIOD / 2;   
        
        -- Second run
        WAIT UNTIL tb_start = '1';
        WAIT FOR CLOCK_PERIOD / 2;
        ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure;
        
        WAIT UNTIL tb_done = '1';
        ASSERT tb_z0 = std_logic_vector(to_unsigned(20, 8))  REPORT "Failed: Z0 was not 0x14"  severity failure;
        ASSERT tb_z1 = std_logic_vector(to_unsigned(400, 8)) REPORT "Failed: Z1 was not 0x190" severity failure;
        ASSERT tb_z2 = std_logic_vector(to_unsigned(0, 8))   REPORT "Failed: Z2 was not 0"     severity failure;
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))   REPORT "Failed: Z3 was not 0"     severity failure;
        WAIT UNTIL tb_done = '0';
        WAIT FOR CLOCK_PERIOD / 2;
        
        -- Thrid run
        WAIT UNTIL tb_start = '1';
        WAIT FOR CLOCK_PERIOD / 2; 
        ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        
        WAIT UNTIL tb_done = '1';
        ASSERT tb_z0 = std_logic_vector(to_unsigned(20, 8))  REPORT "Failed: Z0 was not 0x14"  severity failure;
        ASSERT tb_z1 = std_logic_vector(to_unsigned(400, 8)) REPORT "Failed: Z1 was not 0x190" severity failure;
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))   REPORT "Failed: Z2 was not 0x9"   severity failure;
        ASSERT tb_z3 = std_logic_vector(to_unsigned(0, 8))   REPORT "Failed: Z3 was not 0"     severity failure;
        WAIT UNTIL tb_done = '0';
        WAIT FOR CLOCK_PERIOD / 2;    
        
        -- Fourth run
        WAIT UNTIL tb_start = '1';
        WAIT FOR CLOCK_PERIOD / 2; 
        ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        
        WAIT UNTIL tb_done = '1';
        ASSERT tb_z0 = std_logic_vector(to_unsigned(20, 8))  REPORT "Failed: Z0 was not 0x14"  severity failure;
        ASSERT tb_z1 = std_logic_vector(to_unsigned(400, 8)) REPORT "Failed: Z1 was not 0x190" severity failure;
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))   REPORT "Failed: Z2 was not 0x9"   severity failure;
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "Failed: Z3 was not 0x1A"  severity failure;
        WAIT UNTIL tb_done = '0';
        WAIT FOR CLOCK_PERIOD / 2;    
        
        -- Fifth run
        WAIT UNTIL tb_start = '1';
        WAIT FOR CLOCK_PERIOD / 2; 
        ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
        ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
        ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
        ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
        
        WAIT UNTIL tb_done = '1';
        ASSERT tb_z0 = std_logic_vector(to_unsigned(400, 8)) REPORT "Failed: Z0 was not 0x190" severity failure;
        ASSERT tb_z1 = std_logic_vector(to_unsigned(400, 8)) REPORT "Failed: Z1 was not 0x190" severity failure;
        ASSERT tb_z2 = std_logic_vector(to_unsigned(9, 8))   REPORT "Failed: Z2 was not 0x9"   severity failure;
        ASSERT tb_z3 = std_logic_vector(to_unsigned(26, 8))  REPORT "Failed: Z3 was not 0x1A"  severity failure;
        WAIT UNTIL tb_done = '0';   

        -- FOURTH TEST

         -- First reset
         WAIT UNTIL tb_rst = '1';
         WAIT UNTIL tb_rst = '0';
         ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
         ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
         ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
         ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z3))) severity failure;
         
         -- First run
         WAIT UNTIL tb_start = '1';
         ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
         ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
         ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
         ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure; 
         
         -- Reset after address read
         WAIT UNTIL tb_rst = '1';
         WAIT UNTIL tb_rst = '0';
         ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
         ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
         ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
         ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z3))) severity failure;   
         
         -- Second run
         WAIT UNTIL tb_start = '1';
         ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
         ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
         ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
         ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after the start signal" & integer'image(to_integer(unsigned(tb_z3))) severity failure;
         
         -- Reset at done = '1'
         WAIT UNTIL tb_rst = '1';
         WAIT FOR CLOCK_PERIOD / 2;
         ASSERT tb_z0 = "00000000" REPORT "Failed: Z0 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z0))) severity failure; 
         ASSERT tb_z1 = "00000000" REPORT "Failed: Z1 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z1))) severity failure; 
         ASSERT tb_z2 = "00000000" REPORT "Failed: Z2 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z2))) severity failure; 
         ASSERT tb_z3 = "00000000" REPORT "Failed: Z3 is not zeroed-out after a reset" & integer'image(to_integer(unsigned(tb_z3))) severity failure;
         WAIT UNTIL tb_rst = '0';

        REPORT "Test passed";
        finish;
    END PROCESS testRoutine;

END projecttb;